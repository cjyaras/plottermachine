module mult(a, b, out);
	input [31:0] a, b;
	output [31:0] out;
	
	wire a0b0;
	wire a0b1;
	wire a0b2;
	wire a0b3;
	wire a0b4;
	wire a0b5;
	wire a0b6;
	wire a0b7;
	wire a0b8;
	wire a0b9;
	wire a0b10;
	wire a0b11;
	wire a0b12;
	wire a0b13;
	wire a0b14;
	wire a0b15;
	wire a0b16;
	wire a0b17;
	wire a0b18;
	wire a0b19;
	wire a0b20;
	wire a0b21;
	wire a0b22;
	wire a0b23;
	wire a0b24;
	wire a0b25;
	wire a0b26;
	wire a0b27;
	wire a0b28;
	wire a0b29;
	wire a0b30;
	wire not_a0b31;
	wire a1b0;
	wire a1b1;
	wire a1b2;
	wire a1b3;
	wire a1b4;
	wire a1b5;
	wire a1b6;
	wire a1b7;
	wire a1b8;
	wire a1b9;
	wire a1b10;
	wire a1b11;
	wire a1b12;
	wire a1b13;
	wire a1b14;
	wire a1b15;
	wire a1b16;
	wire a1b17;
	wire a1b18;
	wire a1b19;
	wire a1b20;
	wire a1b21;
	wire a1b22;
	wire a1b23;
	wire a1b24;
	wire a1b25;
	wire a1b26;
	wire a1b27;
	wire a1b28;
	wire a1b29;
	wire a1b30;
	wire not_a1b31;
	wire a2b0;
	wire a2b1;
	wire a2b2;
	wire a2b3;
	wire a2b4;
	wire a2b5;
	wire a2b6;
	wire a2b7;
	wire a2b8;
	wire a2b9;
	wire a2b10;
	wire a2b11;
	wire a2b12;
	wire a2b13;
	wire a2b14;
	wire a2b15;
	wire a2b16;
	wire a2b17;
	wire a2b18;
	wire a2b19;
	wire a2b20;
	wire a2b21;
	wire a2b22;
	wire a2b23;
	wire a2b24;
	wire a2b25;
	wire a2b26;
	wire a2b27;
	wire a2b28;
	wire a2b29;
	wire a2b30;
	wire not_a2b31;
	wire a3b0;
	wire a3b1;
	wire a3b2;
	wire a3b3;
	wire a3b4;
	wire a3b5;
	wire a3b6;
	wire a3b7;
	wire a3b8;
	wire a3b9;
	wire a3b10;
	wire a3b11;
	wire a3b12;
	wire a3b13;
	wire a3b14;
	wire a3b15;
	wire a3b16;
	wire a3b17;
	wire a3b18;
	wire a3b19;
	wire a3b20;
	wire a3b21;
	wire a3b22;
	wire a3b23;
	wire a3b24;
	wire a3b25;
	wire a3b26;
	wire a3b27;
	wire a3b28;
	wire a3b29;
	wire a3b30;
	wire not_a3b31;
	wire a4b0;
	wire a4b1;
	wire a4b2;
	wire a4b3;
	wire a4b4;
	wire a4b5;
	wire a4b6;
	wire a4b7;
	wire a4b8;
	wire a4b9;
	wire a4b10;
	wire a4b11;
	wire a4b12;
	wire a4b13;
	wire a4b14;
	wire a4b15;
	wire a4b16;
	wire a4b17;
	wire a4b18;
	wire a4b19;
	wire a4b20;
	wire a4b21;
	wire a4b22;
	wire a4b23;
	wire a4b24;
	wire a4b25;
	wire a4b26;
	wire a4b27;
	wire a4b28;
	wire a4b29;
	wire a4b30;
	wire not_a4b31;
	wire a5b0;
	wire a5b1;
	wire a5b2;
	wire a5b3;
	wire a5b4;
	wire a5b5;
	wire a5b6;
	wire a5b7;
	wire a5b8;
	wire a5b9;
	wire a5b10;
	wire a5b11;
	wire a5b12;
	wire a5b13;
	wire a5b14;
	wire a5b15;
	wire a5b16;
	wire a5b17;
	wire a5b18;
	wire a5b19;
	wire a5b20;
	wire a5b21;
	wire a5b22;
	wire a5b23;
	wire a5b24;
	wire a5b25;
	wire a5b26;
	wire a5b27;
	wire a5b28;
	wire a5b29;
	wire a5b30;
	wire not_a5b31;
	wire a6b0;
	wire a6b1;
	wire a6b2;
	wire a6b3;
	wire a6b4;
	wire a6b5;
	wire a6b6;
	wire a6b7;
	wire a6b8;
	wire a6b9;
	wire a6b10;
	wire a6b11;
	wire a6b12;
	wire a6b13;
	wire a6b14;
	wire a6b15;
	wire a6b16;
	wire a6b17;
	wire a6b18;
	wire a6b19;
	wire a6b20;
	wire a6b21;
	wire a6b22;
	wire a6b23;
	wire a6b24;
	wire a6b25;
	wire a6b26;
	wire a6b27;
	wire a6b28;
	wire a6b29;
	wire a6b30;
	wire not_a6b31;
	wire a7b0;
	wire a7b1;
	wire a7b2;
	wire a7b3;
	wire a7b4;
	wire a7b5;
	wire a7b6;
	wire a7b7;
	wire a7b8;
	wire a7b9;
	wire a7b10;
	wire a7b11;
	wire a7b12;
	wire a7b13;
	wire a7b14;
	wire a7b15;
	wire a7b16;
	wire a7b17;
	wire a7b18;
	wire a7b19;
	wire a7b20;
	wire a7b21;
	wire a7b22;
	wire a7b23;
	wire a7b24;
	wire a7b25;
	wire a7b26;
	wire a7b27;
	wire a7b28;
	wire a7b29;
	wire a7b30;
	wire not_a7b31;
	wire a8b0;
	wire a8b1;
	wire a8b2;
	wire a8b3;
	wire a8b4;
	wire a8b5;
	wire a8b6;
	wire a8b7;
	wire a8b8;
	wire a8b9;
	wire a8b10;
	wire a8b11;
	wire a8b12;
	wire a8b13;
	wire a8b14;
	wire a8b15;
	wire a8b16;
	wire a8b17;
	wire a8b18;
	wire a8b19;
	wire a8b20;
	wire a8b21;
	wire a8b22;
	wire a8b23;
	wire a8b24;
	wire a8b25;
	wire a8b26;
	wire a8b27;
	wire a8b28;
	wire a8b29;
	wire a8b30;
	wire not_a8b31;
	wire a9b0;
	wire a9b1;
	wire a9b2;
	wire a9b3;
	wire a9b4;
	wire a9b5;
	wire a9b6;
	wire a9b7;
	wire a9b8;
	wire a9b9;
	wire a9b10;
	wire a9b11;
	wire a9b12;
	wire a9b13;
	wire a9b14;
	wire a9b15;
	wire a9b16;
	wire a9b17;
	wire a9b18;
	wire a9b19;
	wire a9b20;
	wire a9b21;
	wire a9b22;
	wire a9b23;
	wire a9b24;
	wire a9b25;
	wire a9b26;
	wire a9b27;
	wire a9b28;
	wire a9b29;
	wire a9b30;
	wire not_a9b31;
	wire a10b0;
	wire a10b1;
	wire a10b2;
	wire a10b3;
	wire a10b4;
	wire a10b5;
	wire a10b6;
	wire a10b7;
	wire a10b8;
	wire a10b9;
	wire a10b10;
	wire a10b11;
	wire a10b12;
	wire a10b13;
	wire a10b14;
	wire a10b15;
	wire a10b16;
	wire a10b17;
	wire a10b18;
	wire a10b19;
	wire a10b20;
	wire a10b21;
	wire a10b22;
	wire a10b23;
	wire a10b24;
	wire a10b25;
	wire a10b26;
	wire a10b27;
	wire a10b28;
	wire a10b29;
	wire a10b30;
	wire not_a10b31;
	wire a11b0;
	wire a11b1;
	wire a11b2;
	wire a11b3;
	wire a11b4;
	wire a11b5;
	wire a11b6;
	wire a11b7;
	wire a11b8;
	wire a11b9;
	wire a11b10;
	wire a11b11;
	wire a11b12;
	wire a11b13;
	wire a11b14;
	wire a11b15;
	wire a11b16;
	wire a11b17;
	wire a11b18;
	wire a11b19;
	wire a11b20;
	wire a11b21;
	wire a11b22;
	wire a11b23;
	wire a11b24;
	wire a11b25;
	wire a11b26;
	wire a11b27;
	wire a11b28;
	wire a11b29;
	wire a11b30;
	wire not_a11b31;
	wire a12b0;
	wire a12b1;
	wire a12b2;
	wire a12b3;
	wire a12b4;
	wire a12b5;
	wire a12b6;
	wire a12b7;
	wire a12b8;
	wire a12b9;
	wire a12b10;
	wire a12b11;
	wire a12b12;
	wire a12b13;
	wire a12b14;
	wire a12b15;
	wire a12b16;
	wire a12b17;
	wire a12b18;
	wire a12b19;
	wire a12b20;
	wire a12b21;
	wire a12b22;
	wire a12b23;
	wire a12b24;
	wire a12b25;
	wire a12b26;
	wire a12b27;
	wire a12b28;
	wire a12b29;
	wire a12b30;
	wire not_a12b31;
	wire a13b0;
	wire a13b1;
	wire a13b2;
	wire a13b3;
	wire a13b4;
	wire a13b5;
	wire a13b6;
	wire a13b7;
	wire a13b8;
	wire a13b9;
	wire a13b10;
	wire a13b11;
	wire a13b12;
	wire a13b13;
	wire a13b14;
	wire a13b15;
	wire a13b16;
	wire a13b17;
	wire a13b18;
	wire a13b19;
	wire a13b20;
	wire a13b21;
	wire a13b22;
	wire a13b23;
	wire a13b24;
	wire a13b25;
	wire a13b26;
	wire a13b27;
	wire a13b28;
	wire a13b29;
	wire a13b30;
	wire not_a13b31;
	wire a14b0;
	wire a14b1;
	wire a14b2;
	wire a14b3;
	wire a14b4;
	wire a14b5;
	wire a14b6;
	wire a14b7;
	wire a14b8;
	wire a14b9;
	wire a14b10;
	wire a14b11;
	wire a14b12;
	wire a14b13;
	wire a14b14;
	wire a14b15;
	wire a14b16;
	wire a14b17;
	wire a14b18;
	wire a14b19;
	wire a14b20;
	wire a14b21;
	wire a14b22;
	wire a14b23;
	wire a14b24;
	wire a14b25;
	wire a14b26;
	wire a14b27;
	wire a14b28;
	wire a14b29;
	wire a14b30;
	wire not_a14b31;
	wire a15b0;
	wire a15b1;
	wire a15b2;
	wire a15b3;
	wire a15b4;
	wire a15b5;
	wire a15b6;
	wire a15b7;
	wire a15b8;
	wire a15b9;
	wire a15b10;
	wire a15b11;
	wire a15b12;
	wire a15b13;
	wire a15b14;
	wire a15b15;
	wire a15b16;
	wire a15b17;
	wire a15b18;
	wire a15b19;
	wire a15b20;
	wire a15b21;
	wire a15b22;
	wire a15b23;
	wire a15b24;
	wire a15b25;
	wire a15b26;
	wire a15b27;
	wire a15b28;
	wire a15b29;
	wire a15b30;
	wire not_a15b31;
	wire a16b0;
	wire a16b1;
	wire a16b2;
	wire a16b3;
	wire a16b4;
	wire a16b5;
	wire a16b6;
	wire a16b7;
	wire a16b8;
	wire a16b9;
	wire a16b10;
	wire a16b11;
	wire a16b12;
	wire a16b13;
	wire a16b14;
	wire a16b15;
	wire a16b16;
	wire a16b17;
	wire a16b18;
	wire a16b19;
	wire a16b20;
	wire a16b21;
	wire a16b22;
	wire a16b23;
	wire a16b24;
	wire a16b25;
	wire a16b26;
	wire a16b27;
	wire a16b28;
	wire a16b29;
	wire a16b30;
	wire not_a16b31;
	wire a17b0;
	wire a17b1;
	wire a17b2;
	wire a17b3;
	wire a17b4;
	wire a17b5;
	wire a17b6;
	wire a17b7;
	wire a17b8;
	wire a17b9;
	wire a17b10;
	wire a17b11;
	wire a17b12;
	wire a17b13;
	wire a17b14;
	wire a17b15;
	wire a17b16;
	wire a17b17;
	wire a17b18;
	wire a17b19;
	wire a17b20;
	wire a17b21;
	wire a17b22;
	wire a17b23;
	wire a17b24;
	wire a17b25;
	wire a17b26;
	wire a17b27;
	wire a17b28;
	wire a17b29;
	wire a17b30;
	wire not_a17b31;
	wire a18b0;
	wire a18b1;
	wire a18b2;
	wire a18b3;
	wire a18b4;
	wire a18b5;
	wire a18b6;
	wire a18b7;
	wire a18b8;
	wire a18b9;
	wire a18b10;
	wire a18b11;
	wire a18b12;
	wire a18b13;
	wire a18b14;
	wire a18b15;
	wire a18b16;
	wire a18b17;
	wire a18b18;
	wire a18b19;
	wire a18b20;
	wire a18b21;
	wire a18b22;
	wire a18b23;
	wire a18b24;
	wire a18b25;
	wire a18b26;
	wire a18b27;
	wire a18b28;
	wire a18b29;
	wire a18b30;
	wire not_a18b31;
	wire a19b0;
	wire a19b1;
	wire a19b2;
	wire a19b3;
	wire a19b4;
	wire a19b5;
	wire a19b6;
	wire a19b7;
	wire a19b8;
	wire a19b9;
	wire a19b10;
	wire a19b11;
	wire a19b12;
	wire a19b13;
	wire a19b14;
	wire a19b15;
	wire a19b16;
	wire a19b17;
	wire a19b18;
	wire a19b19;
	wire a19b20;
	wire a19b21;
	wire a19b22;
	wire a19b23;
	wire a19b24;
	wire a19b25;
	wire a19b26;
	wire a19b27;
	wire a19b28;
	wire a19b29;
	wire a19b30;
	wire not_a19b31;
	wire a20b0;
	wire a20b1;
	wire a20b2;
	wire a20b3;
	wire a20b4;
	wire a20b5;
	wire a20b6;
	wire a20b7;
	wire a20b8;
	wire a20b9;
	wire a20b10;
	wire a20b11;
	wire a20b12;
	wire a20b13;
	wire a20b14;
	wire a20b15;
	wire a20b16;
	wire a20b17;
	wire a20b18;
	wire a20b19;
	wire a20b20;
	wire a20b21;
	wire a20b22;
	wire a20b23;
	wire a20b24;
	wire a20b25;
	wire a20b26;
	wire a20b27;
	wire a20b28;
	wire a20b29;
	wire a20b30;
	wire not_a20b31;
	wire a21b0;
	wire a21b1;
	wire a21b2;
	wire a21b3;
	wire a21b4;
	wire a21b5;
	wire a21b6;
	wire a21b7;
	wire a21b8;
	wire a21b9;
	wire a21b10;
	wire a21b11;
	wire a21b12;
	wire a21b13;
	wire a21b14;
	wire a21b15;
	wire a21b16;
	wire a21b17;
	wire a21b18;
	wire a21b19;
	wire a21b20;
	wire a21b21;
	wire a21b22;
	wire a21b23;
	wire a21b24;
	wire a21b25;
	wire a21b26;
	wire a21b27;
	wire a21b28;
	wire a21b29;
	wire a21b30;
	wire not_a21b31;
	wire a22b0;
	wire a22b1;
	wire a22b2;
	wire a22b3;
	wire a22b4;
	wire a22b5;
	wire a22b6;
	wire a22b7;
	wire a22b8;
	wire a22b9;
	wire a22b10;
	wire a22b11;
	wire a22b12;
	wire a22b13;
	wire a22b14;
	wire a22b15;
	wire a22b16;
	wire a22b17;
	wire a22b18;
	wire a22b19;
	wire a22b20;
	wire a22b21;
	wire a22b22;
	wire a22b23;
	wire a22b24;
	wire a22b25;
	wire a22b26;
	wire a22b27;
	wire a22b28;
	wire a22b29;
	wire a22b30;
	wire not_a22b31;
	wire a23b0;
	wire a23b1;
	wire a23b2;
	wire a23b3;
	wire a23b4;
	wire a23b5;
	wire a23b6;
	wire a23b7;
	wire a23b8;
	wire a23b9;
	wire a23b10;
	wire a23b11;
	wire a23b12;
	wire a23b13;
	wire a23b14;
	wire a23b15;
	wire a23b16;
	wire a23b17;
	wire a23b18;
	wire a23b19;
	wire a23b20;
	wire a23b21;
	wire a23b22;
	wire a23b23;
	wire a23b24;
	wire a23b25;
	wire a23b26;
	wire a23b27;
	wire a23b28;
	wire a23b29;
	wire a23b30;
	wire not_a23b31;
	wire a24b0;
	wire a24b1;
	wire a24b2;
	wire a24b3;
	wire a24b4;
	wire a24b5;
	wire a24b6;
	wire a24b7;
	wire a24b8;
	wire a24b9;
	wire a24b10;
	wire a24b11;
	wire a24b12;
	wire a24b13;
	wire a24b14;
	wire a24b15;
	wire a24b16;
	wire a24b17;
	wire a24b18;
	wire a24b19;
	wire a24b20;
	wire a24b21;
	wire a24b22;
	wire a24b23;
	wire a24b24;
	wire a24b25;
	wire a24b26;
	wire a24b27;
	wire a24b28;
	wire a24b29;
	wire a24b30;
	wire not_a24b31;
	wire a25b0;
	wire a25b1;
	wire a25b2;
	wire a25b3;
	wire a25b4;
	wire a25b5;
	wire a25b6;
	wire a25b7;
	wire a25b8;
	wire a25b9;
	wire a25b10;
	wire a25b11;
	wire a25b12;
	wire a25b13;
	wire a25b14;
	wire a25b15;
	wire a25b16;
	wire a25b17;
	wire a25b18;
	wire a25b19;
	wire a25b20;
	wire a25b21;
	wire a25b22;
	wire a25b23;
	wire a25b24;
	wire a25b25;
	wire a25b26;
	wire a25b27;
	wire a25b28;
	wire a25b29;
	wire a25b30;
	wire not_a25b31;
	wire a26b0;
	wire a26b1;
	wire a26b2;
	wire a26b3;
	wire a26b4;
	wire a26b5;
	wire a26b6;
	wire a26b7;
	wire a26b8;
	wire a26b9;
	wire a26b10;
	wire a26b11;
	wire a26b12;
	wire a26b13;
	wire a26b14;
	wire a26b15;
	wire a26b16;
	wire a26b17;
	wire a26b18;
	wire a26b19;
	wire a26b20;
	wire a26b21;
	wire a26b22;
	wire a26b23;
	wire a26b24;
	wire a26b25;
	wire a26b26;
	wire a26b27;
	wire a26b28;
	wire a26b29;
	wire a26b30;
	wire not_a26b31;
	wire a27b0;
	wire a27b1;
	wire a27b2;
	wire a27b3;
	wire a27b4;
	wire a27b5;
	wire a27b6;
	wire a27b7;
	wire a27b8;
	wire a27b9;
	wire a27b10;
	wire a27b11;
	wire a27b12;
	wire a27b13;
	wire a27b14;
	wire a27b15;
	wire a27b16;
	wire a27b17;
	wire a27b18;
	wire a27b19;
	wire a27b20;
	wire a27b21;
	wire a27b22;
	wire a27b23;
	wire a27b24;
	wire a27b25;
	wire a27b26;
	wire a27b27;
	wire a27b28;
	wire a27b29;
	wire a27b30;
	wire not_a27b31;
	wire a28b0;
	wire a28b1;
	wire a28b2;
	wire a28b3;
	wire a28b4;
	wire a28b5;
	wire a28b6;
	wire a28b7;
	wire a28b8;
	wire a28b9;
	wire a28b10;
	wire a28b11;
	wire a28b12;
	wire a28b13;
	wire a28b14;
	wire a28b15;
	wire a28b16;
	wire a28b17;
	wire a28b18;
	wire a28b19;
	wire a28b20;
	wire a28b21;
	wire a28b22;
	wire a28b23;
	wire a28b24;
	wire a28b25;
	wire a28b26;
	wire a28b27;
	wire a28b28;
	wire a28b29;
	wire a28b30;
	wire not_a28b31;
	wire a29b0;
	wire a29b1;
	wire a29b2;
	wire a29b3;
	wire a29b4;
	wire a29b5;
	wire a29b6;
	wire a29b7;
	wire a29b8;
	wire a29b9;
	wire a29b10;
	wire a29b11;
	wire a29b12;
	wire a29b13;
	wire a29b14;
	wire a29b15;
	wire a29b16;
	wire a29b17;
	wire a29b18;
	wire a29b19;
	wire a29b20;
	wire a29b21;
	wire a29b22;
	wire a29b23;
	wire a29b24;
	wire a29b25;
	wire a29b26;
	wire a29b27;
	wire a29b28;
	wire a29b29;
	wire a29b30;
	wire not_a29b31;
	wire a30b0;
	wire a30b1;
	wire a30b2;
	wire a30b3;
	wire a30b4;
	wire a30b5;
	wire a30b6;
	wire a30b7;
	wire a30b8;
	wire a30b9;
	wire a30b10;
	wire a30b11;
	wire a30b12;
	wire a30b13;
	wire a30b14;
	wire a30b15;
	wire a30b16;
	wire a30b17;
	wire a30b18;
	wire a30b19;
	wire a30b20;
	wire a30b21;
	wire a30b22;
	wire a30b23;
	wire a30b24;
	wire a30b25;
	wire a30b26;
	wire a30b27;
	wire a30b28;
	wire a30b29;
	wire a30b30;
	wire not_a30b31;
	wire not_a31b0;
	wire not_a31b1;
	wire not_a31b2;
	wire not_a31b3;
	wire not_a31b4;
	wire not_a31b5;
	wire not_a31b6;
	wire not_a31b7;
	wire not_a31b8;
	wire not_a31b9;
	wire not_a31b10;
	wire not_a31b11;
	wire not_a31b12;
	wire not_a31b13;
	wire not_a31b14;
	wire not_a31b15;
	wire not_a31b16;
	wire not_a31b17;
	wire not_a31b18;
	wire not_a31b19;
	wire not_a31b20;
	wire not_a31b21;
	wire not_a31b22;
	wire not_a31b23;
	wire not_a31b24;
	wire not_a31b25;
	wire not_a31b26;
	wire not_a31b27;
	wire not_a31b28;
	wire not_a31b29;
	wire not_a31b30;
	wire a31b31;
	wire w_1_1_1;
	wire w_1_2_1;
	wire w_1_2_2;
	wire w_1_3_1;
	wire w_1_3_2;
	wire w_1_4_1;
	wire w_1_4_2;
	wire w_1_5_1;
	wire w_1_4_3;
	wire w_1_5_2;
	wire w_1_5_3;
	wire w_1_6_1;
	wire w_1_5_4;
	wire w_1_6_2;
	wire w_1_6_3;
	wire w_1_7_1;
	wire w_1_6_4;
	wire w_1_7_2;
	wire w_1_7_3;
	wire w_1_8_1;
	wire w_1_7_4;
	wire w_1_8_2;
	wire w_1_7_5;
	wire w_1_8_3;
	wire w_1_8_4;
	wire w_1_9_1;
	wire w_1_8_5;
	wire w_1_9_2;
	wire w_1_8_6;
	wire w_1_9_3;
	wire w_1_9_4;
	wire w_1_10_1;
	wire w_1_9_5;
	wire w_1_10_2;
	wire w_1_9_6;
	wire w_1_10_3;
	wire w_1_10_4;
	wire w_1_11_1;
	wire w_1_10_5;
	wire w_1_11_2;
	wire w_1_10_6;
	wire w_1_11_3;
	wire w_1_10_7;
	wire w_1_11_4;
	wire w_1_11_5;
	wire w_1_12_1;
	wire w_1_11_6;
	wire w_1_12_2;
	wire w_1_11_7;
	wire w_1_12_3;
	wire w_1_11_8;
	wire w_1_12_4;
	wire w_1_12_5;
	wire w_1_13_1;
	wire w_1_12_6;
	wire w_1_13_2;
	wire w_1_12_7;
	wire w_1_13_3;
	wire w_1_12_8;
	wire w_1_13_4;
	wire w_1_13_5;
	wire w_1_14_1;
	wire w_1_13_6;
	wire w_1_14_2;
	wire w_1_13_7;
	wire w_1_14_3;
	wire w_1_13_8;
	wire w_1_14_4;
	wire w_1_13_9;
	wire w_1_14_5;
	wire w_1_14_6;
	wire w_1_15_1;
	wire w_1_14_7;
	wire w_1_15_2;
	wire w_1_14_8;
	wire w_1_15_3;
	wire w_1_14_9;
	wire w_1_15_4;
	wire w_1_14_10;
	wire w_1_15_5;
	wire w_1_15_6;
	wire w_1_16_1;
	wire w_1_15_7;
	wire w_1_16_2;
	wire w_1_15_8;
	wire w_1_16_3;
	wire w_1_15_9;
	wire w_1_16_4;
	wire w_1_15_10;
	wire w_1_16_5;
	wire w_1_16_6;
	wire w_1_17_1;
	wire w_1_16_7;
	wire w_1_17_2;
	wire w_1_16_8;
	wire w_1_17_3;
	wire w_1_16_9;
	wire w_1_17_4;
	wire w_1_16_10;
	wire w_1_17_5;
	wire w_1_16_11;
	wire w_1_17_6;
	wire w_1_17_7;
	wire w_1_18_1;
	wire w_1_17_8;
	wire w_1_18_2;
	wire w_1_17_9;
	wire w_1_18_3;
	wire w_1_17_10;
	wire w_1_18_4;
	wire w_1_17_11;
	wire w_1_18_5;
	wire w_1_17_12;
	wire w_1_18_6;
	wire w_1_18_7;
	wire w_1_19_1;
	wire w_1_18_8;
	wire w_1_19_2;
	wire w_1_18_9;
	wire w_1_19_3;
	wire w_1_18_10;
	wire w_1_19_4;
	wire w_1_18_11;
	wire w_1_19_5;
	wire w_1_18_12;
	wire w_1_19_6;
	wire w_1_19_7;
	wire w_1_20_1;
	wire w_1_19_8;
	wire w_1_20_2;
	wire w_1_19_9;
	wire w_1_20_3;
	wire w_1_19_10;
	wire w_1_20_4;
	wire w_1_19_11;
	wire w_1_20_5;
	wire w_1_19_12;
	wire w_1_20_6;
	wire w_1_19_13;
	wire w_1_20_7;
	wire w_1_20_8;
	wire w_1_21_1;
	wire w_1_20_9;
	wire w_1_21_2;
	wire w_1_20_10;
	wire w_1_21_3;
	wire w_1_20_11;
	wire w_1_21_4;
	wire w_1_20_12;
	wire w_1_21_5;
	wire w_1_20_13;
	wire w_1_21_6;
	wire w_1_20_14;
	wire w_1_21_7;
	wire w_1_21_8;
	wire w_1_22_1;
	wire w_1_21_9;
	wire w_1_22_2;
	wire w_1_21_10;
	wire w_1_22_3;
	wire w_1_21_11;
	wire w_1_22_4;
	wire w_1_21_12;
	wire w_1_22_5;
	wire w_1_21_13;
	wire w_1_22_6;
	wire w_1_21_14;
	wire w_1_22_7;
	wire w_1_22_8;
	wire w_1_23_1;
	wire w_1_22_9;
	wire w_1_23_2;
	wire w_1_22_10;
	wire w_1_23_3;
	wire w_1_22_11;
	wire w_1_23_4;
	wire w_1_22_12;
	wire w_1_23_5;
	wire w_1_22_13;
	wire w_1_23_6;
	wire w_1_22_14;
	wire w_1_23_7;
	wire w_1_22_15;
	wire w_1_23_8;
	wire w_1_23_9;
	wire w_1_24_1;
	wire w_1_23_10;
	wire w_1_24_2;
	wire w_1_23_11;
	wire w_1_24_3;
	wire w_1_23_12;
	wire w_1_24_4;
	wire w_1_23_13;
	wire w_1_24_5;
	wire w_1_23_14;
	wire w_1_24_6;
	wire w_1_23_15;
	wire w_1_24_7;
	wire w_1_23_16;
	wire w_1_24_8;
	wire w_1_24_9;
	wire w_1_25_1;
	wire w_1_24_10;
	wire w_1_25_2;
	wire w_1_24_11;
	wire w_1_25_3;
	wire w_1_24_12;
	wire w_1_25_4;
	wire w_1_24_13;
	wire w_1_25_5;
	wire w_1_24_14;
	wire w_1_25_6;
	wire w_1_24_15;
	wire w_1_25_7;
	wire w_1_24_16;
	wire w_1_25_8;
	wire w_1_25_9;
	wire w_1_26_1;
	wire w_1_25_10;
	wire w_1_26_2;
	wire w_1_25_11;
	wire w_1_26_3;
	wire w_1_25_12;
	wire w_1_26_4;
	wire w_1_25_13;
	wire w_1_26_5;
	wire w_1_25_14;
	wire w_1_26_6;
	wire w_1_25_15;
	wire w_1_26_7;
	wire w_1_25_16;
	wire w_1_26_8;
	wire w_1_25_17;
	wire w_1_26_9;
	wire w_1_26_10;
	wire w_1_27_1;
	wire w_1_26_11;
	wire w_1_27_2;
	wire w_1_26_12;
	wire w_1_27_3;
	wire w_1_26_13;
	wire w_1_27_4;
	wire w_1_26_14;
	wire w_1_27_5;
	wire w_1_26_15;
	wire w_1_27_6;
	wire w_1_26_16;
	wire w_1_27_7;
	wire w_1_26_17;
	wire w_1_27_8;
	wire w_1_26_18;
	wire w_1_27_9;
	wire w_1_27_10;
	wire w_1_28_1;
	wire w_1_27_11;
	wire w_1_28_2;
	wire w_1_27_12;
	wire w_1_28_3;
	wire w_1_27_13;
	wire w_1_28_4;
	wire w_1_27_14;
	wire w_1_28_5;
	wire w_1_27_15;
	wire w_1_28_6;
	wire w_1_27_16;
	wire w_1_28_7;
	wire w_1_27_17;
	wire w_1_28_8;
	wire w_1_27_18;
	wire w_1_28_9;
	wire w_1_28_10;
	wire w_1_29_1;
	wire w_1_28_11;
	wire w_1_29_2;
	wire w_1_28_12;
	wire w_1_29_3;
	wire w_1_28_13;
	wire w_1_29_4;
	wire w_1_28_14;
	wire w_1_29_5;
	wire w_1_28_15;
	wire w_1_29_6;
	wire w_1_28_16;
	wire w_1_29_7;
	wire w_1_28_17;
	wire w_1_29_8;
	wire w_1_28_18;
	wire w_1_29_9;
	wire w_1_28_19;
	wire w_1_29_10;
	wire w_1_29_11;
	wire w_1_30_1;
	wire w_1_29_12;
	wire w_1_30_2;
	wire w_1_29_13;
	wire w_1_30_3;
	wire w_1_29_14;
	wire w_1_30_4;
	wire w_1_29_15;
	wire w_1_30_5;
	wire w_1_29_16;
	wire w_1_30_6;
	wire w_1_29_17;
	wire w_1_30_7;
	wire w_1_29_18;
	wire w_1_30_8;
	wire w_1_29_19;
	wire w_1_30_9;
	wire w_1_29_20;
	wire w_1_30_10;
	wire w_1_30_11;
	wire w_1_31_1;
	wire w_1_30_12;
	wire w_1_31_2;
	wire w_1_30_13;
	wire w_1_31_3;
	wire w_1_30_14;
	wire w_1_31_4;
	wire w_1_30_15;
	wire w_1_31_5;
	wire w_1_30_16;
	wire w_1_31_6;
	wire w_1_30_17;
	wire w_1_31_7;
	wire w_1_30_18;
	wire w_1_31_8;
	wire w_1_30_19;
	wire w_1_31_9;
	wire w_1_30_20;
	wire w_1_31_10;
	wire w_1_31_11;
	wire w_1_32_1;
	wire w_1_31_12;
	wire w_1_32_2;
	wire w_1_31_13;
	wire w_1_32_3;
	wire w_1_31_14;
	wire w_1_32_4;
	wire w_1_31_15;
	wire w_1_32_5;
	wire w_1_31_16;
	wire w_1_32_6;
	wire w_1_31_17;
	wire w_1_32_7;
	wire w_1_31_18;
	wire w_1_32_8;
	wire w_1_31_19;
	wire w_1_32_9;
	wire w_1_31_20;
	wire w_1_32_10;
	wire w_1_31_21;
	wire w_1_32_11;
	wire w_1_32_12;
	wire w_1_33_1;
	wire w_1_32_13;
	wire w_1_33_2;
	wire w_1_32_14;
	wire w_1_33_3;
	wire w_1_32_15;
	wire w_1_33_4;
	wire w_1_32_16;
	wire w_1_33_5;
	wire w_1_32_17;
	wire w_1_33_6;
	wire w_1_32_18;
	wire w_1_33_7;
	wire w_1_32_19;
	wire w_1_33_8;
	wire w_1_32_20;
	wire w_1_33_9;
	wire w_1_32_21;
	wire w_1_33_10;
	wire w_1_32_22;
	wire w_1_33_11;
	wire w_1_33_12;
	wire w_1_34_1;
	wire w_1_33_13;
	wire w_1_34_2;
	wire w_1_33_14;
	wire w_1_34_3;
	wire w_1_33_15;
	wire w_1_34_4;
	wire w_1_33_16;
	wire w_1_34_5;
	wire w_1_33_17;
	wire w_1_34_6;
	wire w_1_33_18;
	wire w_1_34_7;
	wire w_1_33_19;
	wire w_1_34_8;
	wire w_1_33_20;
	wire w_1_34_9;
	wire w_1_33_21;
	wire w_1_34_10;
	wire w_1_34_11;
	wire w_1_35_1;
	wire w_1_34_12;
	wire w_1_35_2;
	wire w_1_34_13;
	wire w_1_35_3;
	wire w_1_34_14;
	wire w_1_35_4;
	wire w_1_34_15;
	wire w_1_35_5;
	wire w_1_34_16;
	wire w_1_35_6;
	wire w_1_34_17;
	wire w_1_35_7;
	wire w_1_34_18;
	wire w_1_35_8;
	wire w_1_34_19;
	wire w_1_35_9;
	wire w_1_34_20;
	wire w_1_35_10;
	wire w_1_35_11;
	wire w_1_36_1;
	wire w_1_35_12;
	wire w_1_36_2;
	wire w_1_35_13;
	wire w_1_36_3;
	wire w_1_35_14;
	wire w_1_36_4;
	wire w_1_35_15;
	wire w_1_36_5;
	wire w_1_35_16;
	wire w_1_36_6;
	wire w_1_35_17;
	wire w_1_36_7;
	wire w_1_35_18;
	wire w_1_36_8;
	wire w_1_35_19;
	wire w_1_36_9;
	wire w_1_36_10;
	wire w_1_37_1;
	wire w_1_36_11;
	wire w_1_37_2;
	wire w_1_36_12;
	wire w_1_37_3;
	wire w_1_36_13;
	wire w_1_37_4;
	wire w_1_36_14;
	wire w_1_37_5;
	wire w_1_36_15;
	wire w_1_37_6;
	wire w_1_36_16;
	wire w_1_37_7;
	wire w_1_36_17;
	wire w_1_37_8;
	wire w_1_36_18;
	wire w_1_37_9;
	wire w_1_37_10;
	wire w_1_38_1;
	wire w_1_37_11;
	wire w_1_38_2;
	wire w_1_37_12;
	wire w_1_38_3;
	wire w_1_37_13;
	wire w_1_38_4;
	wire w_1_37_14;
	wire w_1_38_5;
	wire w_1_37_15;
	wire w_1_38_6;
	wire w_1_37_16;
	wire w_1_38_7;
	wire w_1_37_17;
	wire w_1_38_8;
	wire w_1_37_18;
	wire w_1_38_9;
	wire w_1_38_10;
	wire w_1_39_1;
	wire w_1_38_11;
	wire w_1_39_2;
	wire w_1_38_12;
	wire w_1_39_3;
	wire w_1_38_13;
	wire w_1_39_4;
	wire w_1_38_14;
	wire w_1_39_5;
	wire w_1_38_15;
	wire w_1_39_6;
	wire w_1_38_16;
	wire w_1_39_7;
	wire w_1_38_17;
	wire w_1_39_8;
	wire w_1_39_9;
	wire w_1_40_1;
	wire w_1_39_10;
	wire w_1_40_2;
	wire w_1_39_11;
	wire w_1_40_3;
	wire w_1_39_12;
	wire w_1_40_4;
	wire w_1_39_13;
	wire w_1_40_5;
	wire w_1_39_14;
	wire w_1_40_6;
	wire w_1_39_15;
	wire w_1_40_7;
	wire w_1_39_16;
	wire w_1_40_8;
	wire w_1_40_9;
	wire w_1_41_1;
	wire w_1_40_10;
	wire w_1_41_2;
	wire w_1_40_11;
	wire w_1_41_3;
	wire w_1_40_12;
	wire w_1_41_4;
	wire w_1_40_13;
	wire w_1_41_5;
	wire w_1_40_14;
	wire w_1_41_6;
	wire w_1_40_15;
	wire w_1_41_7;
	wire w_1_40_16;
	wire w_1_41_8;
	wire w_1_41_9;
	wire w_1_42_1;
	wire w_1_41_10;
	wire w_1_42_2;
	wire w_1_41_11;
	wire w_1_42_3;
	wire w_1_41_12;
	wire w_1_42_4;
	wire w_1_41_13;
	wire w_1_42_5;
	wire w_1_41_14;
	wire w_1_42_6;
	wire w_1_41_15;
	wire w_1_42_7;
	wire w_1_42_8;
	wire w_1_43_1;
	wire w_1_42_9;
	wire w_1_43_2;
	wire w_1_42_10;
	wire w_1_43_3;
	wire w_1_42_11;
	wire w_1_43_4;
	wire w_1_42_12;
	wire w_1_43_5;
	wire w_1_42_13;
	wire w_1_43_6;
	wire w_1_42_14;
	wire w_1_43_7;
	wire w_1_43_8;
	wire w_1_44_1;
	wire w_1_43_9;
	wire w_1_44_2;
	wire w_1_43_10;
	wire w_1_44_3;
	wire w_1_43_11;
	wire w_1_44_4;
	wire w_1_43_12;
	wire w_1_44_5;
	wire w_1_43_13;
	wire w_1_44_6;
	wire w_1_43_14;
	wire w_1_44_7;
	wire w_1_44_8;
	wire w_1_45_1;
	wire w_1_44_9;
	wire w_1_45_2;
	wire w_1_44_10;
	wire w_1_45_3;
	wire w_1_44_11;
	wire w_1_45_4;
	wire w_1_44_12;
	wire w_1_45_5;
	wire w_1_44_13;
	wire w_1_45_6;
	wire w_1_45_7;
	wire w_1_46_1;
	wire w_1_45_8;
	wire w_1_46_2;
	wire w_1_45_9;
	wire w_1_46_3;
	wire w_1_45_10;
	wire w_1_46_4;
	wire w_1_45_11;
	wire w_1_46_5;
	wire w_1_45_12;
	wire w_1_46_6;
	wire w_1_46_7;
	wire w_1_47_1;
	wire w_1_46_8;
	wire w_1_47_2;
	wire w_1_46_9;
	wire w_1_47_3;
	wire w_1_46_10;
	wire w_1_47_4;
	wire w_1_46_11;
	wire w_1_47_5;
	wire w_1_46_12;
	wire w_1_47_6;
	wire w_1_47_7;
	wire w_1_48_1;
	wire w_1_47_8;
	wire w_1_48_2;
	wire w_1_47_9;
	wire w_1_48_3;
	wire w_1_47_10;
	wire w_1_48_4;
	wire w_1_47_11;
	wire w_1_48_5;
	wire w_1_48_6;
	wire w_1_49_1;
	wire w_1_48_7;
	wire w_1_49_2;
	wire w_1_48_8;
	wire w_1_49_3;
	wire w_1_48_9;
	wire w_1_49_4;
	wire w_1_48_10;
	wire w_1_49_5;
	wire w_1_49_6;
	wire w_1_50_1;
	wire w_1_49_7;
	wire w_1_50_2;
	wire w_1_49_8;
	wire w_1_50_3;
	wire w_1_49_9;
	wire w_1_50_4;
	wire w_1_49_10;
	wire w_1_50_5;
	wire w_1_50_6;
	wire w_1_51_1;
	wire w_1_50_7;
	wire w_1_51_2;
	wire w_1_50_8;
	wire w_1_51_3;
	wire w_1_50_9;
	wire w_1_51_4;
	wire w_1_51_5;
	wire w_1_52_1;
	wire w_1_51_6;
	wire w_1_52_2;
	wire w_1_51_7;
	wire w_1_52_3;
	wire w_1_51_8;
	wire w_1_52_4;
	wire w_1_52_5;
	wire w_1_53_1;
	wire w_1_52_6;
	wire w_1_53_2;
	wire w_1_52_7;
	wire w_1_53_3;
	wire w_1_52_8;
	wire w_1_53_4;
	wire w_1_53_5;
	wire w_1_54_1;
	wire w_1_53_6;
	wire w_1_54_2;
	wire w_1_53_7;
	wire w_1_54_3;
	wire w_1_54_4;
	wire w_1_55_1;
	wire w_1_54_5;
	wire w_1_55_2;
	wire w_1_54_6;
	wire w_1_55_3;
	wire w_1_55_4;
	wire w_1_56_1;
	wire w_1_55_5;
	wire w_1_56_2;
	wire w_1_55_6;
	wire w_1_56_3;
	wire w_1_56_4;
	wire w_1_57_1;
	wire w_1_56_5;
	wire w_1_57_2;
	wire w_1_57_3;
	wire w_1_58_1;
	wire w_1_57_4;
	wire w_1_58_2;
	wire w_1_58_3;
	wire w_1_59_1;
	wire w_1_58_4;
	wire w_1_59_2;
	wire w_1_59_3;
	wire w_1_60_1;
	wire w_1_60_2;
	wire w_1_61_1;
	wire w_1_61_2;
	wire w_1_62_1;
	wire w_2_2_1;
	wire w_2_3_1;
	wire w_2_3_2;
	wire w_2_4_1;
	wire w_2_4_2;
	wire w_2_5_1;
	wire w_2_5_2;
	wire w_2_6_1;
	wire w_2_6_2;
	wire w_2_7_1;
	wire w_2_6_3;
	wire w_2_7_2;
	wire w_2_7_3;
	wire w_2_8_1;
	wire w_2_7_4;
	wire w_2_8_2;
	wire w_2_8_3;
	wire w_2_9_1;
	wire w_2_8_4;
	wire w_2_9_2;
	wire w_2_9_3;
	wire w_2_10_1;
	wire w_2_9_4;
	wire w_2_10_2;
	wire w_2_10_3;
	wire w_2_11_1;
	wire w_2_10_4;
	wire w_2_11_2;
	wire w_2_11_3;
	wire w_2_12_1;
	wire w_2_11_4;
	wire w_2_12_2;
	wire w_2_11_5;
	wire w_2_12_3;
	wire w_2_12_4;
	wire w_2_13_1;
	wire w_2_12_5;
	wire w_2_13_2;
	wire w_2_12_6;
	wire w_2_13_3;
	wire w_2_13_4;
	wire w_2_14_1;
	wire w_2_13_5;
	wire w_2_14_2;
	wire w_2_13_6;
	wire w_2_14_3;
	wire w_2_14_4;
	wire w_2_15_1;
	wire w_2_14_5;
	wire w_2_15_2;
	wire w_2_14_6;
	wire w_2_15_3;
	wire w_2_15_4;
	wire w_2_16_1;
	wire w_2_15_5;
	wire w_2_16_2;
	wire w_2_15_6;
	wire w_2_16_3;
	wire w_2_15_7;
	wire w_2_16_4;
	wire w_2_16_5;
	wire w_2_17_1;
	wire w_2_16_6;
	wire w_2_17_2;
	wire w_2_16_7;
	wire w_2_17_3;
	wire w_2_16_8;
	wire w_2_17_4;
	wire w_2_17_5;
	wire w_2_18_1;
	wire w_2_17_6;
	wire w_2_18_2;
	wire w_2_17_7;
	wire w_2_18_3;
	wire w_2_17_8;
	wire w_2_18_4;
	wire w_2_18_5;
	wire w_2_19_1;
	wire w_2_18_6;
	wire w_2_19_2;
	wire w_2_18_7;
	wire w_2_19_3;
	wire w_2_18_8;
	wire w_2_19_4;
	wire w_2_19_5;
	wire w_2_20_1;
	wire w_2_19_6;
	wire w_2_20_2;
	wire w_2_19_7;
	wire w_2_20_3;
	wire w_2_19_8;
	wire w_2_20_4;
	wire w_2_20_5;
	wire w_2_21_1;
	wire w_2_20_6;
	wire w_2_21_2;
	wire w_2_20_7;
	wire w_2_21_3;
	wire w_2_20_8;
	wire w_2_21_4;
	wire w_2_20_9;
	wire w_2_21_5;
	wire w_2_21_6;
	wire w_2_22_1;
	wire w_2_21_7;
	wire w_2_22_2;
	wire w_2_21_8;
	wire w_2_22_3;
	wire w_2_21_9;
	wire w_2_22_4;
	wire w_2_21_10;
	wire w_2_22_5;
	wire w_2_22_6;
	wire w_2_23_1;
	wire w_2_22_7;
	wire w_2_23_2;
	wire w_2_22_8;
	wire w_2_23_3;
	wire w_2_22_9;
	wire w_2_23_4;
	wire w_2_22_10;
	wire w_2_23_5;
	wire w_2_23_6;
	wire w_2_24_1;
	wire w_2_23_7;
	wire w_2_24_2;
	wire w_2_23_8;
	wire w_2_24_3;
	wire w_2_23_9;
	wire w_2_24_4;
	wire w_2_23_10;
	wire w_2_24_5;
	wire w_2_24_6;
	wire w_2_25_1;
	wire w_2_24_7;
	wire w_2_25_2;
	wire w_2_24_8;
	wire w_2_25_3;
	wire w_2_24_9;
	wire w_2_25_4;
	wire w_2_24_10;
	wire w_2_25_5;
	wire w_2_24_11;
	wire w_2_25_6;
	wire w_2_25_7;
	wire w_2_26_1;
	wire w_2_25_8;
	wire w_2_26_2;
	wire w_2_25_9;
	wire w_2_26_3;
	wire w_2_25_10;
	wire w_2_26_4;
	wire w_2_25_11;
	wire w_2_26_5;
	wire w_2_25_12;
	wire w_2_26_6;
	wire w_2_26_7;
	wire w_2_27_1;
	wire w_2_26_8;
	wire w_2_27_2;
	wire w_2_26_9;
	wire w_2_27_3;
	wire w_2_26_10;
	wire w_2_27_4;
	wire w_2_26_11;
	wire w_2_27_5;
	wire w_2_26_12;
	wire w_2_27_6;
	wire w_2_27_7;
	wire w_2_28_1;
	wire w_2_27_8;
	wire w_2_28_2;
	wire w_2_27_9;
	wire w_2_28_3;
	wire w_2_27_10;
	wire w_2_28_4;
	wire w_2_27_11;
	wire w_2_28_5;
	wire w_2_27_12;
	wire w_2_28_6;
	wire w_2_28_7;
	wire w_2_29_1;
	wire w_2_28_8;
	wire w_2_29_2;
	wire w_2_28_9;
	wire w_2_29_3;
	wire w_2_28_10;
	wire w_2_29_4;
	wire w_2_28_11;
	wire w_2_29_5;
	wire w_2_28_12;
	wire w_2_29_6;
	wire w_2_29_7;
	wire w_2_30_1;
	wire w_2_29_8;
	wire w_2_30_2;
	wire w_2_29_9;
	wire w_2_30_3;
	wire w_2_29_10;
	wire w_2_30_4;
	wire w_2_29_11;
	wire w_2_30_5;
	wire w_2_29_12;
	wire w_2_30_6;
	wire w_2_29_13;
	wire w_2_30_7;
	wire w_2_30_8;
	wire w_2_31_1;
	wire w_2_30_9;
	wire w_2_31_2;
	wire w_2_30_10;
	wire w_2_31_3;
	wire w_2_30_11;
	wire w_2_31_4;
	wire w_2_30_12;
	wire w_2_31_5;
	wire w_2_30_13;
	wire w_2_31_6;
	wire w_2_30_14;
	wire w_2_31_7;
	wire w_2_31_8;
	wire w_2_32_1;
	wire w_2_31_9;
	wire w_2_32_2;
	wire w_2_31_10;
	wire w_2_32_3;
	wire w_2_31_11;
	wire w_2_32_4;
	wire w_2_31_12;
	wire w_2_32_5;
	wire w_2_31_13;
	wire w_2_32_6;
	wire w_2_31_14;
	wire w_2_32_7;
	wire w_2_32_8;
	wire w_2_33_1;
	wire w_2_32_9;
	wire w_2_33_2;
	wire w_2_32_10;
	wire w_2_33_3;
	wire w_2_32_11;
	wire w_2_33_4;
	wire w_2_32_12;
	wire w_2_33_5;
	wire w_2_32_13;
	wire w_2_33_6;
	wire w_2_32_14;
	wire w_2_33_7;
	wire w_2_33_8;
	wire w_2_34_1;
	wire w_2_33_9;
	wire w_2_34_2;
	wire w_2_33_10;
	wire w_2_34_3;
	wire w_2_33_11;
	wire w_2_34_4;
	wire w_2_33_12;
	wire w_2_34_5;
	wire w_2_33_13;
	wire w_2_34_6;
	wire w_2_33_14;
	wire w_2_34_7;
	wire w_2_34_8;
	wire w_2_35_1;
	wire w_2_34_9;
	wire w_2_35_2;
	wire w_2_34_10;
	wire w_2_35_3;
	wire w_2_34_11;
	wire w_2_35_4;
	wire w_2_34_12;
	wire w_2_35_5;
	wire w_2_34_13;
	wire w_2_35_6;
	wire w_2_34_14;
	wire w_2_35_7;
	wire w_2_35_8;
	wire w_2_36_1;
	wire w_2_35_9;
	wire w_2_36_2;
	wire w_2_35_10;
	wire w_2_36_3;
	wire w_2_35_11;
	wire w_2_36_4;
	wire w_2_35_12;
	wire w_2_36_5;
	wire w_2_35_13;
	wire w_2_36_6;
	wire w_2_35_14;
	wire w_2_36_7;
	wire w_2_36_8;
	wire w_2_37_1;
	wire w_2_36_9;
	wire w_2_37_2;
	wire w_2_36_10;
	wire w_2_37_3;
	wire w_2_36_11;
	wire w_2_37_4;
	wire w_2_36_12;
	wire w_2_37_5;
	wire w_2_36_13;
	wire w_2_37_6;
	wire w_2_37_7;
	wire w_2_38_1;
	wire w_2_37_8;
	wire w_2_38_2;
	wire w_2_37_9;
	wire w_2_38_3;
	wire w_2_37_10;
	wire w_2_38_4;
	wire w_2_37_11;
	wire w_2_38_5;
	wire w_2_37_12;
	wire w_2_38_6;
	wire w_2_38_7;
	wire w_2_39_1;
	wire w_2_38_8;
	wire w_2_39_2;
	wire w_2_38_9;
	wire w_2_39_3;
	wire w_2_38_10;
	wire w_2_39_4;
	wire w_2_38_11;
	wire w_2_39_5;
	wire w_2_38_12;
	wire w_2_39_6;
	wire w_2_39_7;
	wire w_2_40_1;
	wire w_2_39_8;
	wire w_2_40_2;
	wire w_2_39_9;
	wire w_2_40_3;
	wire w_2_39_10;
	wire w_2_40_4;
	wire w_2_39_11;
	wire w_2_40_5;
	wire w_2_40_6;
	wire w_2_41_1;
	wire w_2_40_7;
	wire w_2_41_2;
	wire w_2_40_8;
	wire w_2_41_3;
	wire w_2_40_9;
	wire w_2_41_4;
	wire w_2_40_10;
	wire w_2_41_5;
	wire w_2_41_6;
	wire w_2_42_1;
	wire w_2_41_7;
	wire w_2_42_2;
	wire w_2_41_8;
	wire w_2_42_3;
	wire w_2_41_9;
	wire w_2_42_4;
	wire w_2_41_10;
	wire w_2_42_5;
	wire w_2_42_6;
	wire w_2_43_1;
	wire w_2_42_7;
	wire w_2_43_2;
	wire w_2_42_8;
	wire w_2_43_3;
	wire w_2_42_9;
	wire w_2_43_4;
	wire w_2_42_10;
	wire w_2_43_5;
	wire w_2_43_6;
	wire w_2_44_1;
	wire w_2_43_7;
	wire w_2_44_2;
	wire w_2_43_8;
	wire w_2_44_3;
	wire w_2_43_9;
	wire w_2_44_4;
	wire w_2_43_10;
	wire w_2_44_5;
	wire w_2_44_6;
	wire w_2_45_1;
	wire w_2_44_7;
	wire w_2_45_2;
	wire w_2_44_8;
	wire w_2_45_3;
	wire w_2_44_9;
	wire w_2_45_4;
	wire w_2_44_10;
	wire w_2_45_5;
	wire w_2_45_6;
	wire w_2_46_1;
	wire w_2_45_7;
	wire w_2_46_2;
	wire w_2_45_8;
	wire w_2_46_3;
	wire w_2_45_9;
	wire w_2_46_4;
	wire w_2_46_5;
	wire w_2_47_1;
	wire w_2_46_6;
	wire w_2_47_2;
	wire w_2_46_7;
	wire w_2_47_3;
	wire w_2_46_8;
	wire w_2_47_4;
	wire w_2_47_5;
	wire w_2_48_1;
	wire w_2_47_6;
	wire w_2_48_2;
	wire w_2_47_7;
	wire w_2_48_3;
	wire w_2_47_8;
	wire w_2_48_4;
	wire w_2_48_5;
	wire w_2_49_1;
	wire w_2_48_6;
	wire w_2_49_2;
	wire w_2_48_7;
	wire w_2_49_3;
	wire w_2_49_4;
	wire w_2_50_1;
	wire w_2_49_5;
	wire w_2_50_2;
	wire w_2_49_6;
	wire w_2_50_3;
	wire w_2_50_4;
	wire w_2_51_1;
	wire w_2_50_5;
	wire w_2_51_2;
	wire w_2_50_6;
	wire w_2_51_3;
	wire w_2_51_4;
	wire w_2_52_1;
	wire w_2_51_5;
	wire w_2_52_2;
	wire w_2_51_6;
	wire w_2_52_3;
	wire w_2_52_4;
	wire w_2_53_1;
	wire w_2_52_5;
	wire w_2_53_2;
	wire w_2_52_6;
	wire w_2_53_3;
	wire w_2_53_4;
	wire w_2_54_1;
	wire w_2_53_5;
	wire w_2_54_2;
	wire w_2_53_6;
	wire w_2_54_3;
	wire w_2_54_4;
	wire w_2_55_1;
	wire w_2_54_5;
	wire w_2_55_2;
	wire w_2_55_3;
	wire w_2_56_1;
	wire w_2_55_4;
	wire w_2_56_2;
	wire w_2_56_3;
	wire w_2_57_1;
	wire w_2_56_4;
	wire w_2_57_2;
	wire w_2_57_3;
	wire w_2_58_1;
	wire w_2_58_2;
	wire w_2_59_1;
	wire w_2_59_2;
	wire w_2_60_1;
	wire w_2_60_2;
	wire w_2_61_1;
	wire w_2_61_2;
	wire w_2_62_1;
	wire w_2_62_2;
	wire w_2_63_1;
	wire w_3_3_1;
	wire w_3_4_1;
	wire w_3_4_2;
	wire w_3_5_1;
	wire w_3_5_2;
	wire w_3_6_1;
	wire w_3_6_2;
	wire w_3_7_1;
	wire w_3_7_2;
	wire w_3_8_1;
	wire w_3_8_2;
	wire w_3_9_1;
	wire w_3_9_2;
	wire w_3_10_1;
	wire w_3_9_3;
	wire w_3_10_2;
	wire w_3_10_3;
	wire w_3_11_1;
	wire w_3_10_4;
	wire w_3_11_2;
	wire w_3_11_3;
	wire w_3_12_1;
	wire w_3_11_4;
	wire w_3_12_2;
	wire w_3_12_3;
	wire w_3_13_1;
	wire w_3_12_4;
	wire w_3_13_2;
	wire w_3_13_3;
	wire w_3_14_1;
	wire w_3_13_4;
	wire w_3_14_2;
	wire w_3_14_3;
	wire w_3_15_1;
	wire w_3_14_4;
	wire w_3_15_2;
	wire w_3_15_3;
	wire w_3_16_1;
	wire w_3_15_4;
	wire w_3_16_2;
	wire w_3_16_3;
	wire w_3_17_1;
	wire w_3_16_4;
	wire w_3_17_2;
	wire w_3_16_5;
	wire w_3_17_3;
	wire w_3_17_4;
	wire w_3_18_1;
	wire w_3_17_5;
	wire w_3_18_2;
	wire w_3_17_6;
	wire w_3_18_3;
	wire w_3_18_4;
	wire w_3_19_1;
	wire w_3_18_5;
	wire w_3_19_2;
	wire w_3_18_6;
	wire w_3_19_3;
	wire w_3_19_4;
	wire w_3_20_1;
	wire w_3_19_5;
	wire w_3_20_2;
	wire w_3_19_6;
	wire w_3_20_3;
	wire w_3_20_4;
	wire w_3_21_1;
	wire w_3_20_5;
	wire w_3_21_2;
	wire w_3_20_6;
	wire w_3_21_3;
	wire w_3_21_4;
	wire w_3_22_1;
	wire w_3_21_5;
	wire w_3_22_2;
	wire w_3_21_6;
	wire w_3_22_3;
	wire w_3_22_4;
	wire w_3_23_1;
	wire w_3_22_5;
	wire w_3_23_2;
	wire w_3_22_6;
	wire w_3_23_3;
	wire w_3_23_4;
	wire w_3_24_1;
	wire w_3_23_5;
	wire w_3_24_2;
	wire w_3_23_6;
	wire w_3_24_3;
	wire w_3_23_7;
	wire w_3_24_4;
	wire w_3_24_5;
	wire w_3_25_1;
	wire w_3_24_6;
	wire w_3_25_2;
	wire w_3_24_7;
	wire w_3_25_3;
	wire w_3_24_8;
	wire w_3_25_4;
	wire w_3_25_5;
	wire w_3_26_1;
	wire w_3_25_6;
	wire w_3_26_2;
	wire w_3_25_7;
	wire w_3_26_3;
	wire w_3_25_8;
	wire w_3_26_4;
	wire w_3_26_5;
	wire w_3_27_1;
	wire w_3_26_6;
	wire w_3_27_2;
	wire w_3_26_7;
	wire w_3_27_3;
	wire w_3_26_8;
	wire w_3_27_4;
	wire w_3_27_5;
	wire w_3_28_1;
	wire w_3_27_6;
	wire w_3_28_2;
	wire w_3_27_7;
	wire w_3_28_3;
	wire w_3_27_8;
	wire w_3_28_4;
	wire w_3_28_5;
	wire w_3_29_1;
	wire w_3_28_6;
	wire w_3_29_2;
	wire w_3_28_7;
	wire w_3_29_3;
	wire w_3_28_8;
	wire w_3_29_4;
	wire w_3_29_5;
	wire w_3_30_1;
	wire w_3_29_6;
	wire w_3_30_2;
	wire w_3_29_7;
	wire w_3_30_3;
	wire w_3_29_8;
	wire w_3_30_4;
	wire w_3_30_5;
	wire w_3_31_1;
	wire w_3_30_6;
	wire w_3_31_2;
	wire w_3_30_7;
	wire w_3_31_3;
	wire w_3_30_8;
	wire w_3_31_4;
	wire w_3_30_9;
	wire w_3_31_5;
	wire w_3_31_6;
	wire w_3_32_1;
	wire w_3_31_7;
	wire w_3_32_2;
	wire w_3_31_8;
	wire w_3_32_3;
	wire w_3_31_9;
	wire w_3_32_4;
	wire w_3_31_10;
	wire w_3_32_5;
	wire w_3_32_6;
	wire w_3_33_1;
	wire w_3_32_7;
	wire w_3_33_2;
	wire w_3_32_8;
	wire w_3_33_3;
	wire w_3_32_9;
	wire w_3_33_4;
	wire w_3_32_10;
	wire w_3_33_5;
	wire w_3_33_6;
	wire w_3_34_1;
	wire w_3_33_7;
	wire w_3_34_2;
	wire w_3_33_8;
	wire w_3_34_3;
	wire w_3_33_9;
	wire w_3_34_4;
	wire w_3_33_10;
	wire w_3_34_5;
	wire w_3_34_6;
	wire w_3_35_1;
	wire w_3_34_7;
	wire w_3_35_2;
	wire w_3_34_8;
	wire w_3_35_3;
	wire w_3_34_9;
	wire w_3_35_4;
	wire w_3_34_10;
	wire w_3_35_5;
	wire w_3_35_6;
	wire w_3_36_1;
	wire w_3_35_7;
	wire w_3_36_2;
	wire w_3_35_8;
	wire w_3_36_3;
	wire w_3_35_9;
	wire w_3_36_4;
	wire w_3_35_10;
	wire w_3_36_5;
	wire w_3_36_6;
	wire w_3_37_1;
	wire w_3_36_7;
	wire w_3_37_2;
	wire w_3_36_8;
	wire w_3_37_3;
	wire w_3_36_9;
	wire w_3_37_4;
	wire w_3_37_5;
	wire w_3_38_1;
	wire w_3_37_6;
	wire w_3_38_2;
	wire w_3_37_7;
	wire w_3_38_3;
	wire w_3_37_8;
	wire w_3_38_4;
	wire w_3_38_5;
	wire w_3_39_1;
	wire w_3_38_6;
	wire w_3_39_2;
	wire w_3_38_7;
	wire w_3_39_3;
	wire w_3_38_8;
	wire w_3_39_4;
	wire w_3_39_5;
	wire w_3_40_1;
	wire w_3_39_6;
	wire w_3_40_2;
	wire w_3_39_7;
	wire w_3_40_3;
	wire w_3_39_8;
	wire w_3_40_4;
	wire w_3_40_5;
	wire w_3_41_1;
	wire w_3_40_6;
	wire w_3_41_2;
	wire w_3_40_7;
	wire w_3_41_3;
	wire w_3_40_8;
	wire w_3_41_4;
	wire w_3_41_5;
	wire w_3_42_1;
	wire w_3_41_6;
	wire w_3_42_2;
	wire w_3_41_7;
	wire w_3_42_3;
	wire w_3_41_8;
	wire w_3_42_4;
	wire w_3_42_5;
	wire w_3_43_1;
	wire w_3_42_6;
	wire w_3_43_2;
	wire w_3_42_7;
	wire w_3_43_3;
	wire w_3_43_4;
	wire w_3_44_1;
	wire w_3_43_5;
	wire w_3_44_2;
	wire w_3_43_6;
	wire w_3_44_3;
	wire w_3_44_4;
	wire w_3_45_1;
	wire w_3_44_5;
	wire w_3_45_2;
	wire w_3_44_6;
	wire w_3_45_3;
	wire w_3_45_4;
	wire w_3_46_1;
	wire w_3_45_5;
	wire w_3_46_2;
	wire w_3_45_6;
	wire w_3_46_3;
	wire w_3_46_4;
	wire w_3_47_1;
	wire w_3_46_5;
	wire w_3_47_2;
	wire w_3_46_6;
	wire w_3_47_3;
	wire w_3_47_4;
	wire w_3_48_1;
	wire w_3_47_5;
	wire w_3_48_2;
	wire w_3_47_6;
	wire w_3_48_3;
	wire w_3_48_4;
	wire w_3_49_1;
	wire w_3_48_5;
	wire w_3_49_2;
	wire w_3_48_6;
	wire w_3_49_3;
	wire w_3_49_4;
	wire w_3_50_1;
	wire w_3_49_5;
	wire w_3_50_2;
	wire w_3_50_3;
	wire w_3_51_1;
	wire w_3_50_4;
	wire w_3_51_2;
	wire w_3_51_3;
	wire w_3_52_1;
	wire w_3_51_4;
	wire w_3_52_2;
	wire w_3_52_3;
	wire w_3_53_1;
	wire w_3_52_4;
	wire w_3_53_2;
	wire w_3_53_3;
	wire w_3_54_1;
	wire w_3_53_4;
	wire w_3_54_2;
	wire w_3_54_3;
	wire w_3_55_1;
	wire w_3_54_4;
	wire w_3_55_2;
	wire w_3_55_3;
	wire w_3_56_1;
	wire w_3_56_2;
	wire w_3_57_1;
	wire w_3_57_2;
	wire w_3_58_1;
	wire w_3_58_2;
	wire w_3_59_1;
	wire w_3_59_2;
	wire w_3_60_1;
	wire w_3_60_2;
	wire w_3_61_1;
	wire w_3_61_2;
	wire w_3_62_1;
	wire w_3_62_2;
	wire w_3_63_1;
	wire w_3_63_2;
	wire w_3_64_1;
	wire w_4_4_1;
	wire w_4_5_1;
	wire w_4_5_2;
	wire w_4_6_1;
	wire w_4_6_2;
	wire w_4_7_1;
	wire w_4_7_2;
	wire w_4_8_1;
	wire w_4_8_2;
	wire w_4_9_1;
	wire w_4_9_2;
	wire w_4_10_1;
	wire w_4_10_2;
	wire w_4_11_1;
	wire w_4_11_2;
	wire w_4_12_1;
	wire w_4_12_2;
	wire w_4_13_1;
	wire w_4_13_2;
	wire w_4_14_1;
	wire w_4_14_2;
	wire w_4_15_1;
	wire w_4_14_3;
	wire w_4_15_2;
	wire w_4_15_3;
	wire w_4_16_1;
	wire w_4_15_4;
	wire w_4_16_2;
	wire w_4_16_3;
	wire w_4_17_1;
	wire w_4_16_4;
	wire w_4_17_2;
	wire w_4_17_3;
	wire w_4_18_1;
	wire w_4_17_4;
	wire w_4_18_2;
	wire w_4_18_3;
	wire w_4_19_1;
	wire w_4_18_4;
	wire w_4_19_2;
	wire w_4_19_3;
	wire w_4_20_1;
	wire w_4_19_4;
	wire w_4_20_2;
	wire w_4_20_3;
	wire w_4_21_1;
	wire w_4_20_4;
	wire w_4_21_2;
	wire w_4_21_3;
	wire w_4_22_1;
	wire w_4_21_4;
	wire w_4_22_2;
	wire w_4_22_3;
	wire w_4_23_1;
	wire w_4_22_4;
	wire w_4_23_2;
	wire w_4_23_3;
	wire w_4_24_1;
	wire w_4_23_4;
	wire w_4_24_2;
	wire w_4_24_3;
	wire w_4_25_1;
	wire w_4_24_4;
	wire w_4_25_2;
	wire w_4_24_5;
	wire w_4_25_3;
	wire w_4_25_4;
	wire w_4_26_1;
	wire w_4_25_5;
	wire w_4_26_2;
	wire w_4_25_6;
	wire w_4_26_3;
	wire w_4_26_4;
	wire w_4_27_1;
	wire w_4_26_5;
	wire w_4_27_2;
	wire w_4_26_6;
	wire w_4_27_3;
	wire w_4_27_4;
	wire w_4_28_1;
	wire w_4_27_5;
	wire w_4_28_2;
	wire w_4_27_6;
	wire w_4_28_3;
	wire w_4_28_4;
	wire w_4_29_1;
	wire w_4_28_5;
	wire w_4_29_2;
	wire w_4_28_6;
	wire w_4_29_3;
	wire w_4_29_4;
	wire w_4_30_1;
	wire w_4_29_5;
	wire w_4_30_2;
	wire w_4_29_6;
	wire w_4_30_3;
	wire w_4_30_4;
	wire w_4_31_1;
	wire w_4_30_5;
	wire w_4_31_2;
	wire w_4_30_6;
	wire w_4_31_3;
	wire w_4_31_4;
	wire w_4_32_1;
	wire w_4_31_5;
	wire w_4_32_2;
	wire w_4_31_6;
	wire w_4_32_3;
	wire w_4_32_4;
	wire w_4_33_1;
	wire w_4_32_5;
	wire w_4_33_2;
	wire w_4_32_6;
	wire w_4_33_3;
	wire w_4_33_4;
	wire w_4_34_1;
	wire w_4_33_5;
	wire w_4_34_2;
	wire w_4_33_6;
	wire w_4_34_3;
	wire w_4_34_4;
	wire w_4_35_1;
	wire w_4_34_5;
	wire w_4_35_2;
	wire w_4_34_6;
	wire w_4_35_3;
	wire w_4_35_4;
	wire w_4_36_1;
	wire w_4_35_5;
	wire w_4_36_2;
	wire w_4_35_6;
	wire w_4_36_3;
	wire w_4_36_4;
	wire w_4_37_1;
	wire w_4_36_5;
	wire w_4_37_2;
	wire w_4_36_6;
	wire w_4_37_3;
	wire w_4_37_4;
	wire w_4_38_1;
	wire w_4_37_5;
	wire w_4_38_2;
	wire w_4_37_6;
	wire w_4_38_3;
	wire w_4_38_4;
	wire w_4_39_1;
	wire w_4_38_5;
	wire w_4_39_2;
	wire w_4_38_6;
	wire w_4_39_3;
	wire w_4_39_4;
	wire w_4_40_1;
	wire w_4_39_5;
	wire w_4_40_2;
	wire w_4_39_6;
	wire w_4_40_3;
	wire w_4_40_4;
	wire w_4_41_1;
	wire w_4_40_5;
	wire w_4_41_2;
	wire w_4_40_6;
	wire w_4_41_3;
	wire w_4_41_4;
	wire w_4_42_1;
	wire w_4_41_5;
	wire w_4_42_2;
	wire w_4_41_6;
	wire w_4_42_3;
	wire w_4_42_4;
	wire w_4_43_1;
	wire w_4_42_5;
	wire w_4_43_2;
	wire w_4_42_6;
	wire w_4_43_3;
	wire w_4_43_4;
	wire w_4_44_1;
	wire w_4_43_5;
	wire w_4_44_2;
	wire w_4_44_3;
	wire w_4_45_1;
	wire w_4_44_4;
	wire w_4_45_2;
	wire w_4_45_3;
	wire w_4_46_1;
	wire w_4_45_4;
	wire w_4_46_2;
	wire w_4_46_3;
	wire w_4_47_1;
	wire w_4_46_4;
	wire w_4_47_2;
	wire w_4_47_3;
	wire w_4_48_1;
	wire w_4_47_4;
	wire w_4_48_2;
	wire w_4_48_3;
	wire w_4_49_1;
	wire w_4_48_4;
	wire w_4_49_2;
	wire w_4_49_3;
	wire w_4_50_1;
	wire w_4_49_4;
	wire w_4_50_2;
	wire w_4_50_3;
	wire w_4_51_1;
	wire w_4_50_4;
	wire w_4_51_2;
	wire w_4_51_3;
	wire w_4_52_1;
	wire w_4_52_2;
	wire w_4_53_1;
	wire w_4_53_2;
	wire w_4_54_1;
	wire w_4_54_2;
	wire w_4_55_1;
	wire w_4_55_2;
	wire w_4_56_1;
	wire w_4_56_2;
	wire w_4_57_1;
	wire w_4_57_2;
	wire w_4_58_1;
	wire w_4_58_2;
	wire w_4_59_1;
	wire w_4_59_2;
	wire w_4_60_1;
	wire w_4_60_2;
	wire w_4_61_1;
	wire w_4_61_2;
	wire w_4_62_1;
	wire w_4_62_2;
	wire w_4_63_1;
	wire w_4_63_2;
	wire w_4_64_1;
	wire w_5_5_1;
	wire w_5_6_1;
	wire w_5_6_2;
	wire w_5_7_1;
	wire w_5_7_2;
	wire w_5_8_1;
	wire w_5_8_2;
	wire w_5_9_1;
	wire w_5_9_2;
	wire w_5_10_1;
	wire w_5_10_2;
	wire w_5_11_1;
	wire w_5_11_2;
	wire w_5_12_1;
	wire w_5_12_2;
	wire w_5_13_1;
	wire w_5_13_2;
	wire w_5_14_1;
	wire w_5_14_2;
	wire w_5_15_1;
	wire w_5_15_2;
	wire w_5_16_1;
	wire w_5_16_2;
	wire w_5_17_1;
	wire w_5_17_2;
	wire w_5_18_1;
	wire w_5_18_2;
	wire w_5_19_1;
	wire w_5_19_2;
	wire w_5_20_1;
	wire w_5_20_2;
	wire w_5_21_1;
	wire w_5_21_2;
	wire w_5_22_1;
	wire w_5_21_3;
	wire w_5_22_2;
	wire w_5_22_3;
	wire w_5_23_1;
	wire w_5_22_4;
	wire w_5_23_2;
	wire w_5_23_3;
	wire w_5_24_1;
	wire w_5_23_4;
	wire w_5_24_2;
	wire w_5_24_3;
	wire w_5_25_1;
	wire w_5_24_4;
	wire w_5_25_2;
	wire w_5_25_3;
	wire w_5_26_1;
	wire w_5_25_4;
	wire w_5_26_2;
	wire w_5_26_3;
	wire w_5_27_1;
	wire w_5_26_4;
	wire w_5_27_2;
	wire w_5_27_3;
	wire w_5_28_1;
	wire w_5_27_4;
	wire w_5_28_2;
	wire w_5_28_3;
	wire w_5_29_1;
	wire w_5_28_4;
	wire w_5_29_2;
	wire w_5_29_3;
	wire w_5_30_1;
	wire w_5_29_4;
	wire w_5_30_2;
	wire w_5_30_3;
	wire w_5_31_1;
	wire w_5_30_4;
	wire w_5_31_2;
	wire w_5_31_3;
	wire w_5_32_1;
	wire w_5_31_4;
	wire w_5_32_2;
	wire w_5_32_3;
	wire w_5_33_1;
	wire w_5_32_4;
	wire w_5_33_2;
	wire w_5_33_3;
	wire w_5_34_1;
	wire w_5_33_4;
	wire w_5_34_2;
	wire w_5_34_3;
	wire w_5_35_1;
	wire w_5_34_4;
	wire w_5_35_2;
	wire w_5_35_3;
	wire w_5_36_1;
	wire w_5_35_4;
	wire w_5_36_2;
	wire w_5_36_3;
	wire w_5_37_1;
	wire w_5_36_4;
	wire w_5_37_2;
	wire w_5_37_3;
	wire w_5_38_1;
	wire w_5_37_4;
	wire w_5_38_2;
	wire w_5_38_3;
	wire w_5_39_1;
	wire w_5_38_4;
	wire w_5_39_2;
	wire w_5_39_3;
	wire w_5_40_1;
	wire w_5_39_4;
	wire w_5_40_2;
	wire w_5_40_3;
	wire w_5_41_1;
	wire w_5_40_4;
	wire w_5_41_2;
	wire w_5_41_3;
	wire w_5_42_1;
	wire w_5_41_4;
	wire w_5_42_2;
	wire w_5_42_3;
	wire w_5_43_1;
	wire w_5_42_4;
	wire w_5_43_2;
	wire w_5_43_3;
	wire w_5_44_1;
	wire w_5_43_4;
	wire w_5_44_2;
	wire w_5_44_3;
	wire w_5_45_1;
	wire w_5_44_4;
	wire w_5_45_2;
	wire w_5_45_3;
	wire w_5_46_1;
	wire w_5_46_2;
	wire w_5_47_1;
	wire w_5_47_2;
	wire w_5_48_1;
	wire w_5_48_2;
	wire w_5_49_1;
	wire w_5_49_2;
	wire w_5_50_1;
	wire w_5_50_2;
	wire w_5_51_1;
	wire w_5_51_2;
	wire w_5_52_1;
	wire w_5_52_2;
	wire w_5_53_1;
	wire w_5_53_2;
	wire w_5_54_1;
	wire w_5_54_2;
	wire w_5_55_1;
	wire w_5_55_2;
	wire w_5_56_1;
	wire w_5_56_2;
	wire w_5_57_1;
	wire w_5_57_2;
	wire w_5_58_1;
	wire w_5_58_2;
	wire w_5_59_1;
	wire w_5_59_2;
	wire w_5_60_1;
	wire w_5_60_2;
	wire w_5_61_1;
	wire w_5_61_2;
	wire w_5_62_1;
	wire w_5_62_2;
	wire w_5_63_1;
	wire w_5_63_2;
	wire w_5_64_1;
	wire w_5_64_2;
	wire w_5_65_1;
	wire w_6_6_1;
	wire w_6_7_1;
	wire w_6_7_2;
	wire w_6_8_1;
	wire w_6_8_2;
	wire w_6_9_1;
	wire w_6_9_2;
	wire w_6_10_1;
	wire w_6_10_2;
	wire w_6_11_1;
	wire w_6_11_2;
	wire w_6_12_1;
	wire w_6_12_2;
	wire w_6_13_1;
	wire w_6_13_2;
	wire w_6_14_1;
	wire w_6_14_2;
	wire w_6_15_1;
	wire w_6_15_2;
	wire w_6_16_1;
	wire w_6_16_2;
	wire w_6_17_1;
	wire w_6_17_2;
	wire w_6_18_1;
	wire w_6_18_2;
	wire w_6_19_1;
	wire w_6_19_2;
	wire w_6_20_1;
	wire w_6_20_2;
	wire w_6_21_1;
	wire w_6_21_2;
	wire w_6_22_1;
	wire w_6_22_2;
	wire w_6_23_1;
	wire w_6_23_2;
	wire w_6_24_1;
	wire w_6_24_2;
	wire w_6_25_1;
	wire w_6_25_2;
	wire w_6_26_1;
	wire w_6_26_2;
	wire w_6_27_1;
	wire w_6_27_2;
	wire w_6_28_1;
	wire w_6_28_2;
	wire w_6_29_1;
	wire w_6_29_2;
	wire w_6_30_1;
	wire w_6_30_2;
	wire w_6_31_1;
	wire w_6_31_2;
	wire w_6_32_1;
	wire w_6_31_3;
	wire w_6_32_2;
	wire w_6_32_3;
	wire w_6_33_1;
	wire w_6_32_4;
	wire w_6_33_2;
	wire w_6_33_3;
	wire w_6_34_1;
	wire w_6_33_4;
	wire w_6_34_2;
	wire w_6_34_3;
	wire w_6_35_1;
	wire w_6_34_4;
	wire w_6_35_2;
	wire w_6_35_3;
	wire w_6_36_1;
	wire w_6_35_4;
	wire w_6_36_2;
	wire w_6_36_3;
	wire w_6_37_1;
	wire w_6_36_4;
	wire w_6_37_2;
	wire w_6_37_3;
	wire w_6_38_1;
	wire w_6_38_2;
	wire w_6_39_1;
	wire w_6_39_2;
	wire w_6_40_1;
	wire w_6_40_2;
	wire w_6_41_1;
	wire w_6_41_2;
	wire w_6_42_1;
	wire w_6_42_2;
	wire w_6_43_1;
	wire w_6_43_2;
	wire w_6_44_1;
	wire w_6_44_2;
	wire w_6_45_1;
	wire w_6_45_2;
	wire w_6_46_1;
	wire w_6_46_2;
	wire w_6_47_1;
	wire w_6_47_2;
	wire w_6_48_1;
	wire w_6_48_2;
	wire w_6_49_1;
	wire w_6_49_2;
	wire w_6_50_1;
	wire w_6_50_2;
	wire w_6_51_1;
	wire w_6_51_2;
	wire w_6_52_1;
	wire w_6_52_2;
	wire w_6_53_1;
	wire w_6_53_2;
	wire w_6_54_1;
	wire w_6_54_2;
	wire w_6_55_1;
	wire w_6_55_2;
	wire w_6_56_1;
	wire w_6_56_2;
	wire w_6_57_1;
	wire w_6_57_2;
	wire w_6_58_1;
	wire w_6_58_2;
	wire w_6_59_1;
	wire w_6_59_2;
	wire w_6_60_1;
	wire w_6_60_2;
	wire w_6_61_1;
	wire w_6_61_2;
	wire w_6_62_1;
	wire w_6_62_2;
	wire w_6_63_1;
	wire w_6_63_2;
	wire w_6_64_1;
	wire w_6_64_2;
	wire w_6_65_1;
	wire w_7_7_1;
	wire w_7_8_1;
	wire w_7_8_2;
	wire w_7_9_1;
	wire w_7_9_2;
	wire w_7_10_1;
	wire w_7_10_2;
	wire w_7_11_1;
	wire w_7_11_2;
	wire w_7_12_1;
	wire w_7_12_2;
	wire w_7_13_1;
	wire w_7_13_2;
	wire w_7_14_1;
	wire w_7_14_2;
	wire w_7_15_1;
	wire w_7_15_2;
	wire w_7_16_1;
	wire w_7_16_2;
	wire w_7_17_1;
	wire w_7_17_2;
	wire w_7_18_1;
	wire w_7_18_2;
	wire w_7_19_1;
	wire w_7_19_2;
	wire w_7_20_1;
	wire w_7_20_2;
	wire w_7_21_1;
	wire w_7_21_2;
	wire w_7_22_1;
	wire w_7_22_2;
	wire w_7_23_1;
	wire w_7_23_2;
	wire w_7_24_1;
	wire w_7_24_2;
	wire w_7_25_1;
	wire w_7_25_2;
	wire w_7_26_1;
	wire w_7_26_2;
	wire w_7_27_1;
	wire w_7_27_2;
	wire w_7_28_1;
	wire w_7_28_2;
	wire w_7_29_1;
	wire w_7_29_2;
	wire w_7_30_1;
	wire w_7_30_2;
	wire w_7_31_1;
	wire w_7_31_2;
	wire w_7_32_1;
	wire w_7_32_2;
	wire w_7_33_1;
	wire w_7_33_2;
	wire w_7_34_1;
	wire w_7_34_2;
	wire w_7_35_1;
	wire w_7_35_2;
	wire w_7_36_1;
	wire w_7_36_2;
	wire w_7_37_1;
	wire w_7_37_2;
	wire w_7_38_1;
	wire w_7_38_2;
	wire w_7_39_1;
	wire w_7_39_2;
	wire w_7_40_1;
	wire w_7_40_2;
	wire w_7_41_1;
	wire w_7_41_2;
	wire w_7_42_1;
	wire w_7_42_2;
	wire w_7_43_1;
	wire w_7_43_2;
	wire w_7_44_1;
	wire w_7_44_2;
	wire w_7_45_1;
	wire w_7_45_2;
	wire w_7_46_1;
	wire w_7_46_2;
	wire w_7_47_1;
	wire w_7_47_2;
	wire w_7_48_1;
	wire w_7_48_2;
	wire w_7_49_1;
	wire w_7_49_2;
	wire w_7_50_1;
	wire w_7_50_2;
	wire w_7_51_1;
	wire w_7_51_2;
	wire w_7_52_1;
	wire w_7_52_2;
	wire w_7_53_1;
	wire w_7_53_2;
	wire w_7_54_1;
	wire w_7_54_2;
	wire w_7_55_1;
	wire w_7_55_2;
	wire w_7_56_1;
	wire w_7_56_2;
	wire w_7_57_1;
	wire w_7_57_2;
	wire w_7_58_1;
	wire w_7_58_2;
	wire w_7_59_1;
	wire w_7_59_2;
	wire w_7_60_1;
	wire w_7_60_2;
	wire w_7_61_1;
	wire w_7_61_2;
	wire w_7_62_1;
	wire w_7_62_2;
	wire w_7_63_1;
	wire w_7_63_2;
	wire w_7_64_1;
	wire w_7_64_2;
	wire w_7_65_1;
	wire w_7_65_2;
	wire w_7_66_1;
	wire w_8_8_1;
	wire w_8_9_1;
	wire w_8_9_2;
	wire w_8_10_1;
	wire w_8_10_2;
	wire w_8_11_1;
	wire w_8_11_2;
	wire w_8_12_1;
	wire w_8_12_2;
	wire w_8_13_1;
	wire w_8_13_2;
	wire w_8_14_1;
	wire w_8_14_2;
	wire w_8_15_1;
	wire w_8_15_2;
	wire w_8_16_1;
	wire w_8_16_2;
	wire w_8_17_1;
	wire w_8_17_2;
	wire w_8_18_1;
	wire w_8_18_2;
	wire w_8_19_1;
	wire w_8_19_2;
	wire w_8_20_1;
	wire w_8_20_2;
	wire w_8_21_1;
	wire w_8_21_2;
	wire w_8_22_1;
	wire w_8_22_2;
	wire w_8_23_1;
	wire w_8_23_2;
	wire w_8_24_1;
	wire w_8_24_2;
	wire w_8_25_1;
	wire w_8_25_2;
	wire w_8_26_1;
	wire w_8_26_2;
	wire w_8_27_1;
	wire w_8_27_2;
	wire w_8_28_1;
	wire w_8_28_2;
	wire w_8_29_1;
	wire w_8_29_2;
	wire w_8_30_1;
	wire w_8_30_2;
	wire w_8_31_1;
	wire w_8_31_2;
	wire w_8_32_1;
	wire w_8_32_2;
	wire w_8_33_1;
	wire w_8_33_2;
	wire w_8_34_1;
	wire w_8_34_2;
	wire w_8_35_1;
	wire w_8_35_2;
	wire w_8_36_1;
	wire w_8_36_2;
	wire w_8_37_1;
	wire w_8_37_2;
	wire w_8_38_1;
	wire w_8_38_2;
	wire w_8_39_1;
	wire w_8_39_2;
	wire w_8_40_1;
	wire w_8_40_2;
	wire w_8_41_1;
	wire w_8_41_2;
	wire w_8_42_1;
	wire w_8_42_2;
	wire w_8_43_1;
	wire w_8_43_2;
	wire w_8_44_1;
	wire w_8_44_2;
	wire w_8_45_1;
	wire w_8_45_2;
	wire w_8_46_1;
	wire w_8_46_2;
	wire w_8_47_1;
	wire w_8_47_2;
	wire w_8_48_1;
	wire w_8_48_2;
	wire w_8_49_1;
	wire w_8_49_2;
	wire w_8_50_1;
	wire w_8_50_2;
	wire w_8_51_1;
	wire w_8_51_2;
	wire w_8_52_1;
	wire w_8_52_2;
	wire w_8_53_1;
	wire w_8_53_2;
	wire w_8_54_1;
	wire w_8_54_2;
	wire w_8_55_1;
	wire w_8_55_2;
	wire w_8_56_1;
	wire w_8_56_2;
	wire w_8_57_1;
	wire w_8_57_2;
	wire w_8_58_1;
	wire w_8_58_2;
	wire w_8_59_1;
	wire w_8_59_2;
	wire w_8_60_1;
	wire w_8_60_2;
	wire w_8_61_1;
	wire w_8_61_2;
	wire w_8_62_1;
	wire w_8_62_2;
	wire w_8_63_1;
	wire w_8_63_2;
	wire w_8_64_1;
	wire w_8_64_2;
	wire w_8_65_1;
	wire w_8_65_2;
	wire w_8_66_1;
	wire [63:0] result1, result2;

	and and_a0b0(a0b0, a[0], b[0]);
	and and_a0b1(a0b1, a[0], b[1]);
	and and_a0b2(a0b2, a[0], b[2]);
	and and_a0b3(a0b3, a[0], b[3]);
	and and_a0b4(a0b4, a[0], b[4]);
	and and_a0b5(a0b5, a[0], b[5]);
	and and_a0b6(a0b6, a[0], b[6]);
	and and_a0b7(a0b7, a[0], b[7]);
	and and_a0b8(a0b8, a[0], b[8]);
	and and_a0b9(a0b9, a[0], b[9]);
	and and_a0b10(a0b10, a[0], b[10]);
	and and_a0b11(a0b11, a[0], b[11]);
	and and_a0b12(a0b12, a[0], b[12]);
	and and_a0b13(a0b13, a[0], b[13]);
	and and_a0b14(a0b14, a[0], b[14]);
	and and_a0b15(a0b15, a[0], b[15]);
	and and_a0b16(a0b16, a[0], b[16]);
	and and_a0b17(a0b17, a[0], b[17]);
	and and_a0b18(a0b18, a[0], b[18]);
	and and_a0b19(a0b19, a[0], b[19]);
	and and_a0b20(a0b20, a[0], b[20]);
	and and_a0b21(a0b21, a[0], b[21]);
	and and_a0b22(a0b22, a[0], b[22]);
	and and_a0b23(a0b23, a[0], b[23]);
	and and_a0b24(a0b24, a[0], b[24]);
	and and_a0b25(a0b25, a[0], b[25]);
	and and_a0b26(a0b26, a[0], b[26]);
	and and_a0b27(a0b27, a[0], b[27]);
	and and_a0b28(a0b28, a[0], b[28]);
	and and_a0b29(a0b29, a[0], b[29]);
	and and_a0b30(a0b30, a[0], b[30]);
	nand nand_a0b31(not_a0b31, a[0], b[31]);
	and and_a1b0(a1b0, a[1], b[0]);
	and and_a1b1(a1b1, a[1], b[1]);
	and and_a1b2(a1b2, a[1], b[2]);
	and and_a1b3(a1b3, a[1], b[3]);
	and and_a1b4(a1b4, a[1], b[4]);
	and and_a1b5(a1b5, a[1], b[5]);
	and and_a1b6(a1b6, a[1], b[6]);
	and and_a1b7(a1b7, a[1], b[7]);
	and and_a1b8(a1b8, a[1], b[8]);
	and and_a1b9(a1b9, a[1], b[9]);
	and and_a1b10(a1b10, a[1], b[10]);
	and and_a1b11(a1b11, a[1], b[11]);
	and and_a1b12(a1b12, a[1], b[12]);
	and and_a1b13(a1b13, a[1], b[13]);
	and and_a1b14(a1b14, a[1], b[14]);
	and and_a1b15(a1b15, a[1], b[15]);
	and and_a1b16(a1b16, a[1], b[16]);
	and and_a1b17(a1b17, a[1], b[17]);
	and and_a1b18(a1b18, a[1], b[18]);
	and and_a1b19(a1b19, a[1], b[19]);
	and and_a1b20(a1b20, a[1], b[20]);
	and and_a1b21(a1b21, a[1], b[21]);
	and and_a1b22(a1b22, a[1], b[22]);
	and and_a1b23(a1b23, a[1], b[23]);
	and and_a1b24(a1b24, a[1], b[24]);
	and and_a1b25(a1b25, a[1], b[25]);
	and and_a1b26(a1b26, a[1], b[26]);
	and and_a1b27(a1b27, a[1], b[27]);
	and and_a1b28(a1b28, a[1], b[28]);
	and and_a1b29(a1b29, a[1], b[29]);
	and and_a1b30(a1b30, a[1], b[30]);
	nand nand_a1b31(not_a1b31, a[1], b[31]);
	and and_a2b0(a2b0, a[2], b[0]);
	and and_a2b1(a2b1, a[2], b[1]);
	and and_a2b2(a2b2, a[2], b[2]);
	and and_a2b3(a2b3, a[2], b[3]);
	and and_a2b4(a2b4, a[2], b[4]);
	and and_a2b5(a2b5, a[2], b[5]);
	and and_a2b6(a2b6, a[2], b[6]);
	and and_a2b7(a2b7, a[2], b[7]);
	and and_a2b8(a2b8, a[2], b[8]);
	and and_a2b9(a2b9, a[2], b[9]);
	and and_a2b10(a2b10, a[2], b[10]);
	and and_a2b11(a2b11, a[2], b[11]);
	and and_a2b12(a2b12, a[2], b[12]);
	and and_a2b13(a2b13, a[2], b[13]);
	and and_a2b14(a2b14, a[2], b[14]);
	and and_a2b15(a2b15, a[2], b[15]);
	and and_a2b16(a2b16, a[2], b[16]);
	and and_a2b17(a2b17, a[2], b[17]);
	and and_a2b18(a2b18, a[2], b[18]);
	and and_a2b19(a2b19, a[2], b[19]);
	and and_a2b20(a2b20, a[2], b[20]);
	and and_a2b21(a2b21, a[2], b[21]);
	and and_a2b22(a2b22, a[2], b[22]);
	and and_a2b23(a2b23, a[2], b[23]);
	and and_a2b24(a2b24, a[2], b[24]);
	and and_a2b25(a2b25, a[2], b[25]);
	and and_a2b26(a2b26, a[2], b[26]);
	and and_a2b27(a2b27, a[2], b[27]);
	and and_a2b28(a2b28, a[2], b[28]);
	and and_a2b29(a2b29, a[2], b[29]);
	and and_a2b30(a2b30, a[2], b[30]);
	nand nand_a2b31(not_a2b31, a[2], b[31]);
	and and_a3b0(a3b0, a[3], b[0]);
	and and_a3b1(a3b1, a[3], b[1]);
	and and_a3b2(a3b2, a[3], b[2]);
	and and_a3b3(a3b3, a[3], b[3]);
	and and_a3b4(a3b4, a[3], b[4]);
	and and_a3b5(a3b5, a[3], b[5]);
	and and_a3b6(a3b6, a[3], b[6]);
	and and_a3b7(a3b7, a[3], b[7]);
	and and_a3b8(a3b8, a[3], b[8]);
	and and_a3b9(a3b9, a[3], b[9]);
	and and_a3b10(a3b10, a[3], b[10]);
	and and_a3b11(a3b11, a[3], b[11]);
	and and_a3b12(a3b12, a[3], b[12]);
	and and_a3b13(a3b13, a[3], b[13]);
	and and_a3b14(a3b14, a[3], b[14]);
	and and_a3b15(a3b15, a[3], b[15]);
	and and_a3b16(a3b16, a[3], b[16]);
	and and_a3b17(a3b17, a[3], b[17]);
	and and_a3b18(a3b18, a[3], b[18]);
	and and_a3b19(a3b19, a[3], b[19]);
	and and_a3b20(a3b20, a[3], b[20]);
	and and_a3b21(a3b21, a[3], b[21]);
	and and_a3b22(a3b22, a[3], b[22]);
	and and_a3b23(a3b23, a[3], b[23]);
	and and_a3b24(a3b24, a[3], b[24]);
	and and_a3b25(a3b25, a[3], b[25]);
	and and_a3b26(a3b26, a[3], b[26]);
	and and_a3b27(a3b27, a[3], b[27]);
	and and_a3b28(a3b28, a[3], b[28]);
	and and_a3b29(a3b29, a[3], b[29]);
	and and_a3b30(a3b30, a[3], b[30]);
	nand nand_a3b31(not_a3b31, a[3], b[31]);
	and and_a4b0(a4b0, a[4], b[0]);
	and and_a4b1(a4b1, a[4], b[1]);
	and and_a4b2(a4b2, a[4], b[2]);
	and and_a4b3(a4b3, a[4], b[3]);
	and and_a4b4(a4b4, a[4], b[4]);
	and and_a4b5(a4b5, a[4], b[5]);
	and and_a4b6(a4b6, a[4], b[6]);
	and and_a4b7(a4b7, a[4], b[7]);
	and and_a4b8(a4b8, a[4], b[8]);
	and and_a4b9(a4b9, a[4], b[9]);
	and and_a4b10(a4b10, a[4], b[10]);
	and and_a4b11(a4b11, a[4], b[11]);
	and and_a4b12(a4b12, a[4], b[12]);
	and and_a4b13(a4b13, a[4], b[13]);
	and and_a4b14(a4b14, a[4], b[14]);
	and and_a4b15(a4b15, a[4], b[15]);
	and and_a4b16(a4b16, a[4], b[16]);
	and and_a4b17(a4b17, a[4], b[17]);
	and and_a4b18(a4b18, a[4], b[18]);
	and and_a4b19(a4b19, a[4], b[19]);
	and and_a4b20(a4b20, a[4], b[20]);
	and and_a4b21(a4b21, a[4], b[21]);
	and and_a4b22(a4b22, a[4], b[22]);
	and and_a4b23(a4b23, a[4], b[23]);
	and and_a4b24(a4b24, a[4], b[24]);
	and and_a4b25(a4b25, a[4], b[25]);
	and and_a4b26(a4b26, a[4], b[26]);
	and and_a4b27(a4b27, a[4], b[27]);
	and and_a4b28(a4b28, a[4], b[28]);
	and and_a4b29(a4b29, a[4], b[29]);
	and and_a4b30(a4b30, a[4], b[30]);
	nand nand_a4b31(not_a4b31, a[4], b[31]);
	and and_a5b0(a5b0, a[5], b[0]);
	and and_a5b1(a5b1, a[5], b[1]);
	and and_a5b2(a5b2, a[5], b[2]);
	and and_a5b3(a5b3, a[5], b[3]);
	and and_a5b4(a5b4, a[5], b[4]);
	and and_a5b5(a5b5, a[5], b[5]);
	and and_a5b6(a5b6, a[5], b[6]);
	and and_a5b7(a5b7, a[5], b[7]);
	and and_a5b8(a5b8, a[5], b[8]);
	and and_a5b9(a5b9, a[5], b[9]);
	and and_a5b10(a5b10, a[5], b[10]);
	and and_a5b11(a5b11, a[5], b[11]);
	and and_a5b12(a5b12, a[5], b[12]);
	and and_a5b13(a5b13, a[5], b[13]);
	and and_a5b14(a5b14, a[5], b[14]);
	and and_a5b15(a5b15, a[5], b[15]);
	and and_a5b16(a5b16, a[5], b[16]);
	and and_a5b17(a5b17, a[5], b[17]);
	and and_a5b18(a5b18, a[5], b[18]);
	and and_a5b19(a5b19, a[5], b[19]);
	and and_a5b20(a5b20, a[5], b[20]);
	and and_a5b21(a5b21, a[5], b[21]);
	and and_a5b22(a5b22, a[5], b[22]);
	and and_a5b23(a5b23, a[5], b[23]);
	and and_a5b24(a5b24, a[5], b[24]);
	and and_a5b25(a5b25, a[5], b[25]);
	and and_a5b26(a5b26, a[5], b[26]);
	and and_a5b27(a5b27, a[5], b[27]);
	and and_a5b28(a5b28, a[5], b[28]);
	and and_a5b29(a5b29, a[5], b[29]);
	and and_a5b30(a5b30, a[5], b[30]);
	nand nand_a5b31(not_a5b31, a[5], b[31]);
	and and_a6b0(a6b0, a[6], b[0]);
	and and_a6b1(a6b1, a[6], b[1]);
	and and_a6b2(a6b2, a[6], b[2]);
	and and_a6b3(a6b3, a[6], b[3]);
	and and_a6b4(a6b4, a[6], b[4]);
	and and_a6b5(a6b5, a[6], b[5]);
	and and_a6b6(a6b6, a[6], b[6]);
	and and_a6b7(a6b7, a[6], b[7]);
	and and_a6b8(a6b8, a[6], b[8]);
	and and_a6b9(a6b9, a[6], b[9]);
	and and_a6b10(a6b10, a[6], b[10]);
	and and_a6b11(a6b11, a[6], b[11]);
	and and_a6b12(a6b12, a[6], b[12]);
	and and_a6b13(a6b13, a[6], b[13]);
	and and_a6b14(a6b14, a[6], b[14]);
	and and_a6b15(a6b15, a[6], b[15]);
	and and_a6b16(a6b16, a[6], b[16]);
	and and_a6b17(a6b17, a[6], b[17]);
	and and_a6b18(a6b18, a[6], b[18]);
	and and_a6b19(a6b19, a[6], b[19]);
	and and_a6b20(a6b20, a[6], b[20]);
	and and_a6b21(a6b21, a[6], b[21]);
	and and_a6b22(a6b22, a[6], b[22]);
	and and_a6b23(a6b23, a[6], b[23]);
	and and_a6b24(a6b24, a[6], b[24]);
	and and_a6b25(a6b25, a[6], b[25]);
	and and_a6b26(a6b26, a[6], b[26]);
	and and_a6b27(a6b27, a[6], b[27]);
	and and_a6b28(a6b28, a[6], b[28]);
	and and_a6b29(a6b29, a[6], b[29]);
	and and_a6b30(a6b30, a[6], b[30]);
	nand nand_a6b31(not_a6b31, a[6], b[31]);
	and and_a7b0(a7b0, a[7], b[0]);
	and and_a7b1(a7b1, a[7], b[1]);
	and and_a7b2(a7b2, a[7], b[2]);
	and and_a7b3(a7b3, a[7], b[3]);
	and and_a7b4(a7b4, a[7], b[4]);
	and and_a7b5(a7b5, a[7], b[5]);
	and and_a7b6(a7b6, a[7], b[6]);
	and and_a7b7(a7b7, a[7], b[7]);
	and and_a7b8(a7b8, a[7], b[8]);
	and and_a7b9(a7b9, a[7], b[9]);
	and and_a7b10(a7b10, a[7], b[10]);
	and and_a7b11(a7b11, a[7], b[11]);
	and and_a7b12(a7b12, a[7], b[12]);
	and and_a7b13(a7b13, a[7], b[13]);
	and and_a7b14(a7b14, a[7], b[14]);
	and and_a7b15(a7b15, a[7], b[15]);
	and and_a7b16(a7b16, a[7], b[16]);
	and and_a7b17(a7b17, a[7], b[17]);
	and and_a7b18(a7b18, a[7], b[18]);
	and and_a7b19(a7b19, a[7], b[19]);
	and and_a7b20(a7b20, a[7], b[20]);
	and and_a7b21(a7b21, a[7], b[21]);
	and and_a7b22(a7b22, a[7], b[22]);
	and and_a7b23(a7b23, a[7], b[23]);
	and and_a7b24(a7b24, a[7], b[24]);
	and and_a7b25(a7b25, a[7], b[25]);
	and and_a7b26(a7b26, a[7], b[26]);
	and and_a7b27(a7b27, a[7], b[27]);
	and and_a7b28(a7b28, a[7], b[28]);
	and and_a7b29(a7b29, a[7], b[29]);
	and and_a7b30(a7b30, a[7], b[30]);
	nand nand_a7b31(not_a7b31, a[7], b[31]);
	and and_a8b0(a8b0, a[8], b[0]);
	and and_a8b1(a8b1, a[8], b[1]);
	and and_a8b2(a8b2, a[8], b[2]);
	and and_a8b3(a8b3, a[8], b[3]);
	and and_a8b4(a8b4, a[8], b[4]);
	and and_a8b5(a8b5, a[8], b[5]);
	and and_a8b6(a8b6, a[8], b[6]);
	and and_a8b7(a8b7, a[8], b[7]);
	and and_a8b8(a8b8, a[8], b[8]);
	and and_a8b9(a8b9, a[8], b[9]);
	and and_a8b10(a8b10, a[8], b[10]);
	and and_a8b11(a8b11, a[8], b[11]);
	and and_a8b12(a8b12, a[8], b[12]);
	and and_a8b13(a8b13, a[8], b[13]);
	and and_a8b14(a8b14, a[8], b[14]);
	and and_a8b15(a8b15, a[8], b[15]);
	and and_a8b16(a8b16, a[8], b[16]);
	and and_a8b17(a8b17, a[8], b[17]);
	and and_a8b18(a8b18, a[8], b[18]);
	and and_a8b19(a8b19, a[8], b[19]);
	and and_a8b20(a8b20, a[8], b[20]);
	and and_a8b21(a8b21, a[8], b[21]);
	and and_a8b22(a8b22, a[8], b[22]);
	and and_a8b23(a8b23, a[8], b[23]);
	and and_a8b24(a8b24, a[8], b[24]);
	and and_a8b25(a8b25, a[8], b[25]);
	and and_a8b26(a8b26, a[8], b[26]);
	and and_a8b27(a8b27, a[8], b[27]);
	and and_a8b28(a8b28, a[8], b[28]);
	and and_a8b29(a8b29, a[8], b[29]);
	and and_a8b30(a8b30, a[8], b[30]);
	nand nand_a8b31(not_a8b31, a[8], b[31]);
	and and_a9b0(a9b0, a[9], b[0]);
	and and_a9b1(a9b1, a[9], b[1]);
	and and_a9b2(a9b2, a[9], b[2]);
	and and_a9b3(a9b3, a[9], b[3]);
	and and_a9b4(a9b4, a[9], b[4]);
	and and_a9b5(a9b5, a[9], b[5]);
	and and_a9b6(a9b6, a[9], b[6]);
	and and_a9b7(a9b7, a[9], b[7]);
	and and_a9b8(a9b8, a[9], b[8]);
	and and_a9b9(a9b9, a[9], b[9]);
	and and_a9b10(a9b10, a[9], b[10]);
	and and_a9b11(a9b11, a[9], b[11]);
	and and_a9b12(a9b12, a[9], b[12]);
	and and_a9b13(a9b13, a[9], b[13]);
	and and_a9b14(a9b14, a[9], b[14]);
	and and_a9b15(a9b15, a[9], b[15]);
	and and_a9b16(a9b16, a[9], b[16]);
	and and_a9b17(a9b17, a[9], b[17]);
	and and_a9b18(a9b18, a[9], b[18]);
	and and_a9b19(a9b19, a[9], b[19]);
	and and_a9b20(a9b20, a[9], b[20]);
	and and_a9b21(a9b21, a[9], b[21]);
	and and_a9b22(a9b22, a[9], b[22]);
	and and_a9b23(a9b23, a[9], b[23]);
	and and_a9b24(a9b24, a[9], b[24]);
	and and_a9b25(a9b25, a[9], b[25]);
	and and_a9b26(a9b26, a[9], b[26]);
	and and_a9b27(a9b27, a[9], b[27]);
	and and_a9b28(a9b28, a[9], b[28]);
	and and_a9b29(a9b29, a[9], b[29]);
	and and_a9b30(a9b30, a[9], b[30]);
	nand nand_a9b31(not_a9b31, a[9], b[31]);
	and and_a10b0(a10b0, a[10], b[0]);
	and and_a10b1(a10b1, a[10], b[1]);
	and and_a10b2(a10b2, a[10], b[2]);
	and and_a10b3(a10b3, a[10], b[3]);
	and and_a10b4(a10b4, a[10], b[4]);
	and and_a10b5(a10b5, a[10], b[5]);
	and and_a10b6(a10b6, a[10], b[6]);
	and and_a10b7(a10b7, a[10], b[7]);
	and and_a10b8(a10b8, a[10], b[8]);
	and and_a10b9(a10b9, a[10], b[9]);
	and and_a10b10(a10b10, a[10], b[10]);
	and and_a10b11(a10b11, a[10], b[11]);
	and and_a10b12(a10b12, a[10], b[12]);
	and and_a10b13(a10b13, a[10], b[13]);
	and and_a10b14(a10b14, a[10], b[14]);
	and and_a10b15(a10b15, a[10], b[15]);
	and and_a10b16(a10b16, a[10], b[16]);
	and and_a10b17(a10b17, a[10], b[17]);
	and and_a10b18(a10b18, a[10], b[18]);
	and and_a10b19(a10b19, a[10], b[19]);
	and and_a10b20(a10b20, a[10], b[20]);
	and and_a10b21(a10b21, a[10], b[21]);
	and and_a10b22(a10b22, a[10], b[22]);
	and and_a10b23(a10b23, a[10], b[23]);
	and and_a10b24(a10b24, a[10], b[24]);
	and and_a10b25(a10b25, a[10], b[25]);
	and and_a10b26(a10b26, a[10], b[26]);
	and and_a10b27(a10b27, a[10], b[27]);
	and and_a10b28(a10b28, a[10], b[28]);
	and and_a10b29(a10b29, a[10], b[29]);
	and and_a10b30(a10b30, a[10], b[30]);
	nand nand_a10b31(not_a10b31, a[10], b[31]);
	and and_a11b0(a11b0, a[11], b[0]);
	and and_a11b1(a11b1, a[11], b[1]);
	and and_a11b2(a11b2, a[11], b[2]);
	and and_a11b3(a11b3, a[11], b[3]);
	and and_a11b4(a11b4, a[11], b[4]);
	and and_a11b5(a11b5, a[11], b[5]);
	and and_a11b6(a11b6, a[11], b[6]);
	and and_a11b7(a11b7, a[11], b[7]);
	and and_a11b8(a11b8, a[11], b[8]);
	and and_a11b9(a11b9, a[11], b[9]);
	and and_a11b10(a11b10, a[11], b[10]);
	and and_a11b11(a11b11, a[11], b[11]);
	and and_a11b12(a11b12, a[11], b[12]);
	and and_a11b13(a11b13, a[11], b[13]);
	and and_a11b14(a11b14, a[11], b[14]);
	and and_a11b15(a11b15, a[11], b[15]);
	and and_a11b16(a11b16, a[11], b[16]);
	and and_a11b17(a11b17, a[11], b[17]);
	and and_a11b18(a11b18, a[11], b[18]);
	and and_a11b19(a11b19, a[11], b[19]);
	and and_a11b20(a11b20, a[11], b[20]);
	and and_a11b21(a11b21, a[11], b[21]);
	and and_a11b22(a11b22, a[11], b[22]);
	and and_a11b23(a11b23, a[11], b[23]);
	and and_a11b24(a11b24, a[11], b[24]);
	and and_a11b25(a11b25, a[11], b[25]);
	and and_a11b26(a11b26, a[11], b[26]);
	and and_a11b27(a11b27, a[11], b[27]);
	and and_a11b28(a11b28, a[11], b[28]);
	and and_a11b29(a11b29, a[11], b[29]);
	and and_a11b30(a11b30, a[11], b[30]);
	nand nand_a11b31(not_a11b31, a[11], b[31]);
	and and_a12b0(a12b0, a[12], b[0]);
	and and_a12b1(a12b1, a[12], b[1]);
	and and_a12b2(a12b2, a[12], b[2]);
	and and_a12b3(a12b3, a[12], b[3]);
	and and_a12b4(a12b4, a[12], b[4]);
	and and_a12b5(a12b5, a[12], b[5]);
	and and_a12b6(a12b6, a[12], b[6]);
	and and_a12b7(a12b7, a[12], b[7]);
	and and_a12b8(a12b8, a[12], b[8]);
	and and_a12b9(a12b9, a[12], b[9]);
	and and_a12b10(a12b10, a[12], b[10]);
	and and_a12b11(a12b11, a[12], b[11]);
	and and_a12b12(a12b12, a[12], b[12]);
	and and_a12b13(a12b13, a[12], b[13]);
	and and_a12b14(a12b14, a[12], b[14]);
	and and_a12b15(a12b15, a[12], b[15]);
	and and_a12b16(a12b16, a[12], b[16]);
	and and_a12b17(a12b17, a[12], b[17]);
	and and_a12b18(a12b18, a[12], b[18]);
	and and_a12b19(a12b19, a[12], b[19]);
	and and_a12b20(a12b20, a[12], b[20]);
	and and_a12b21(a12b21, a[12], b[21]);
	and and_a12b22(a12b22, a[12], b[22]);
	and and_a12b23(a12b23, a[12], b[23]);
	and and_a12b24(a12b24, a[12], b[24]);
	and and_a12b25(a12b25, a[12], b[25]);
	and and_a12b26(a12b26, a[12], b[26]);
	and and_a12b27(a12b27, a[12], b[27]);
	and and_a12b28(a12b28, a[12], b[28]);
	and and_a12b29(a12b29, a[12], b[29]);
	and and_a12b30(a12b30, a[12], b[30]);
	nand nand_a12b31(not_a12b31, a[12], b[31]);
	and and_a13b0(a13b0, a[13], b[0]);
	and and_a13b1(a13b1, a[13], b[1]);
	and and_a13b2(a13b2, a[13], b[2]);
	and and_a13b3(a13b3, a[13], b[3]);
	and and_a13b4(a13b4, a[13], b[4]);
	and and_a13b5(a13b5, a[13], b[5]);
	and and_a13b6(a13b6, a[13], b[6]);
	and and_a13b7(a13b7, a[13], b[7]);
	and and_a13b8(a13b8, a[13], b[8]);
	and and_a13b9(a13b9, a[13], b[9]);
	and and_a13b10(a13b10, a[13], b[10]);
	and and_a13b11(a13b11, a[13], b[11]);
	and and_a13b12(a13b12, a[13], b[12]);
	and and_a13b13(a13b13, a[13], b[13]);
	and and_a13b14(a13b14, a[13], b[14]);
	and and_a13b15(a13b15, a[13], b[15]);
	and and_a13b16(a13b16, a[13], b[16]);
	and and_a13b17(a13b17, a[13], b[17]);
	and and_a13b18(a13b18, a[13], b[18]);
	and and_a13b19(a13b19, a[13], b[19]);
	and and_a13b20(a13b20, a[13], b[20]);
	and and_a13b21(a13b21, a[13], b[21]);
	and and_a13b22(a13b22, a[13], b[22]);
	and and_a13b23(a13b23, a[13], b[23]);
	and and_a13b24(a13b24, a[13], b[24]);
	and and_a13b25(a13b25, a[13], b[25]);
	and and_a13b26(a13b26, a[13], b[26]);
	and and_a13b27(a13b27, a[13], b[27]);
	and and_a13b28(a13b28, a[13], b[28]);
	and and_a13b29(a13b29, a[13], b[29]);
	and and_a13b30(a13b30, a[13], b[30]);
	nand nand_a13b31(not_a13b31, a[13], b[31]);
	and and_a14b0(a14b0, a[14], b[0]);
	and and_a14b1(a14b1, a[14], b[1]);
	and and_a14b2(a14b2, a[14], b[2]);
	and and_a14b3(a14b3, a[14], b[3]);
	and and_a14b4(a14b4, a[14], b[4]);
	and and_a14b5(a14b5, a[14], b[5]);
	and and_a14b6(a14b6, a[14], b[6]);
	and and_a14b7(a14b7, a[14], b[7]);
	and and_a14b8(a14b8, a[14], b[8]);
	and and_a14b9(a14b9, a[14], b[9]);
	and and_a14b10(a14b10, a[14], b[10]);
	and and_a14b11(a14b11, a[14], b[11]);
	and and_a14b12(a14b12, a[14], b[12]);
	and and_a14b13(a14b13, a[14], b[13]);
	and and_a14b14(a14b14, a[14], b[14]);
	and and_a14b15(a14b15, a[14], b[15]);
	and and_a14b16(a14b16, a[14], b[16]);
	and and_a14b17(a14b17, a[14], b[17]);
	and and_a14b18(a14b18, a[14], b[18]);
	and and_a14b19(a14b19, a[14], b[19]);
	and and_a14b20(a14b20, a[14], b[20]);
	and and_a14b21(a14b21, a[14], b[21]);
	and and_a14b22(a14b22, a[14], b[22]);
	and and_a14b23(a14b23, a[14], b[23]);
	and and_a14b24(a14b24, a[14], b[24]);
	and and_a14b25(a14b25, a[14], b[25]);
	and and_a14b26(a14b26, a[14], b[26]);
	and and_a14b27(a14b27, a[14], b[27]);
	and and_a14b28(a14b28, a[14], b[28]);
	and and_a14b29(a14b29, a[14], b[29]);
	and and_a14b30(a14b30, a[14], b[30]);
	nand nand_a14b31(not_a14b31, a[14], b[31]);
	and and_a15b0(a15b0, a[15], b[0]);
	and and_a15b1(a15b1, a[15], b[1]);
	and and_a15b2(a15b2, a[15], b[2]);
	and and_a15b3(a15b3, a[15], b[3]);
	and and_a15b4(a15b4, a[15], b[4]);
	and and_a15b5(a15b5, a[15], b[5]);
	and and_a15b6(a15b6, a[15], b[6]);
	and and_a15b7(a15b7, a[15], b[7]);
	and and_a15b8(a15b8, a[15], b[8]);
	and and_a15b9(a15b9, a[15], b[9]);
	and and_a15b10(a15b10, a[15], b[10]);
	and and_a15b11(a15b11, a[15], b[11]);
	and and_a15b12(a15b12, a[15], b[12]);
	and and_a15b13(a15b13, a[15], b[13]);
	and and_a15b14(a15b14, a[15], b[14]);
	and and_a15b15(a15b15, a[15], b[15]);
	and and_a15b16(a15b16, a[15], b[16]);
	and and_a15b17(a15b17, a[15], b[17]);
	and and_a15b18(a15b18, a[15], b[18]);
	and and_a15b19(a15b19, a[15], b[19]);
	and and_a15b20(a15b20, a[15], b[20]);
	and and_a15b21(a15b21, a[15], b[21]);
	and and_a15b22(a15b22, a[15], b[22]);
	and and_a15b23(a15b23, a[15], b[23]);
	and and_a15b24(a15b24, a[15], b[24]);
	and and_a15b25(a15b25, a[15], b[25]);
	and and_a15b26(a15b26, a[15], b[26]);
	and and_a15b27(a15b27, a[15], b[27]);
	and and_a15b28(a15b28, a[15], b[28]);
	and and_a15b29(a15b29, a[15], b[29]);
	and and_a15b30(a15b30, a[15], b[30]);
	nand nand_a15b31(not_a15b31, a[15], b[31]);
	and and_a16b0(a16b0, a[16], b[0]);
	and and_a16b1(a16b1, a[16], b[1]);
	and and_a16b2(a16b2, a[16], b[2]);
	and and_a16b3(a16b3, a[16], b[3]);
	and and_a16b4(a16b4, a[16], b[4]);
	and and_a16b5(a16b5, a[16], b[5]);
	and and_a16b6(a16b6, a[16], b[6]);
	and and_a16b7(a16b7, a[16], b[7]);
	and and_a16b8(a16b8, a[16], b[8]);
	and and_a16b9(a16b9, a[16], b[9]);
	and and_a16b10(a16b10, a[16], b[10]);
	and and_a16b11(a16b11, a[16], b[11]);
	and and_a16b12(a16b12, a[16], b[12]);
	and and_a16b13(a16b13, a[16], b[13]);
	and and_a16b14(a16b14, a[16], b[14]);
	and and_a16b15(a16b15, a[16], b[15]);
	and and_a16b16(a16b16, a[16], b[16]);
	and and_a16b17(a16b17, a[16], b[17]);
	and and_a16b18(a16b18, a[16], b[18]);
	and and_a16b19(a16b19, a[16], b[19]);
	and and_a16b20(a16b20, a[16], b[20]);
	and and_a16b21(a16b21, a[16], b[21]);
	and and_a16b22(a16b22, a[16], b[22]);
	and and_a16b23(a16b23, a[16], b[23]);
	and and_a16b24(a16b24, a[16], b[24]);
	and and_a16b25(a16b25, a[16], b[25]);
	and and_a16b26(a16b26, a[16], b[26]);
	and and_a16b27(a16b27, a[16], b[27]);
	and and_a16b28(a16b28, a[16], b[28]);
	and and_a16b29(a16b29, a[16], b[29]);
	and and_a16b30(a16b30, a[16], b[30]);
	nand nand_a16b31(not_a16b31, a[16], b[31]);
	and and_a17b0(a17b0, a[17], b[0]);
	and and_a17b1(a17b1, a[17], b[1]);
	and and_a17b2(a17b2, a[17], b[2]);
	and and_a17b3(a17b3, a[17], b[3]);
	and and_a17b4(a17b4, a[17], b[4]);
	and and_a17b5(a17b5, a[17], b[5]);
	and and_a17b6(a17b6, a[17], b[6]);
	and and_a17b7(a17b7, a[17], b[7]);
	and and_a17b8(a17b8, a[17], b[8]);
	and and_a17b9(a17b9, a[17], b[9]);
	and and_a17b10(a17b10, a[17], b[10]);
	and and_a17b11(a17b11, a[17], b[11]);
	and and_a17b12(a17b12, a[17], b[12]);
	and and_a17b13(a17b13, a[17], b[13]);
	and and_a17b14(a17b14, a[17], b[14]);
	and and_a17b15(a17b15, a[17], b[15]);
	and and_a17b16(a17b16, a[17], b[16]);
	and and_a17b17(a17b17, a[17], b[17]);
	and and_a17b18(a17b18, a[17], b[18]);
	and and_a17b19(a17b19, a[17], b[19]);
	and and_a17b20(a17b20, a[17], b[20]);
	and and_a17b21(a17b21, a[17], b[21]);
	and and_a17b22(a17b22, a[17], b[22]);
	and and_a17b23(a17b23, a[17], b[23]);
	and and_a17b24(a17b24, a[17], b[24]);
	and and_a17b25(a17b25, a[17], b[25]);
	and and_a17b26(a17b26, a[17], b[26]);
	and and_a17b27(a17b27, a[17], b[27]);
	and and_a17b28(a17b28, a[17], b[28]);
	and and_a17b29(a17b29, a[17], b[29]);
	and and_a17b30(a17b30, a[17], b[30]);
	nand nand_a17b31(not_a17b31, a[17], b[31]);
	and and_a18b0(a18b0, a[18], b[0]);
	and and_a18b1(a18b1, a[18], b[1]);
	and and_a18b2(a18b2, a[18], b[2]);
	and and_a18b3(a18b3, a[18], b[3]);
	and and_a18b4(a18b4, a[18], b[4]);
	and and_a18b5(a18b5, a[18], b[5]);
	and and_a18b6(a18b6, a[18], b[6]);
	and and_a18b7(a18b7, a[18], b[7]);
	and and_a18b8(a18b8, a[18], b[8]);
	and and_a18b9(a18b9, a[18], b[9]);
	and and_a18b10(a18b10, a[18], b[10]);
	and and_a18b11(a18b11, a[18], b[11]);
	and and_a18b12(a18b12, a[18], b[12]);
	and and_a18b13(a18b13, a[18], b[13]);
	and and_a18b14(a18b14, a[18], b[14]);
	and and_a18b15(a18b15, a[18], b[15]);
	and and_a18b16(a18b16, a[18], b[16]);
	and and_a18b17(a18b17, a[18], b[17]);
	and and_a18b18(a18b18, a[18], b[18]);
	and and_a18b19(a18b19, a[18], b[19]);
	and and_a18b20(a18b20, a[18], b[20]);
	and and_a18b21(a18b21, a[18], b[21]);
	and and_a18b22(a18b22, a[18], b[22]);
	and and_a18b23(a18b23, a[18], b[23]);
	and and_a18b24(a18b24, a[18], b[24]);
	and and_a18b25(a18b25, a[18], b[25]);
	and and_a18b26(a18b26, a[18], b[26]);
	and and_a18b27(a18b27, a[18], b[27]);
	and and_a18b28(a18b28, a[18], b[28]);
	and and_a18b29(a18b29, a[18], b[29]);
	and and_a18b30(a18b30, a[18], b[30]);
	nand nand_a18b31(not_a18b31, a[18], b[31]);
	and and_a19b0(a19b0, a[19], b[0]);
	and and_a19b1(a19b1, a[19], b[1]);
	and and_a19b2(a19b2, a[19], b[2]);
	and and_a19b3(a19b3, a[19], b[3]);
	and and_a19b4(a19b4, a[19], b[4]);
	and and_a19b5(a19b5, a[19], b[5]);
	and and_a19b6(a19b6, a[19], b[6]);
	and and_a19b7(a19b7, a[19], b[7]);
	and and_a19b8(a19b8, a[19], b[8]);
	and and_a19b9(a19b9, a[19], b[9]);
	and and_a19b10(a19b10, a[19], b[10]);
	and and_a19b11(a19b11, a[19], b[11]);
	and and_a19b12(a19b12, a[19], b[12]);
	and and_a19b13(a19b13, a[19], b[13]);
	and and_a19b14(a19b14, a[19], b[14]);
	and and_a19b15(a19b15, a[19], b[15]);
	and and_a19b16(a19b16, a[19], b[16]);
	and and_a19b17(a19b17, a[19], b[17]);
	and and_a19b18(a19b18, a[19], b[18]);
	and and_a19b19(a19b19, a[19], b[19]);
	and and_a19b20(a19b20, a[19], b[20]);
	and and_a19b21(a19b21, a[19], b[21]);
	and and_a19b22(a19b22, a[19], b[22]);
	and and_a19b23(a19b23, a[19], b[23]);
	and and_a19b24(a19b24, a[19], b[24]);
	and and_a19b25(a19b25, a[19], b[25]);
	and and_a19b26(a19b26, a[19], b[26]);
	and and_a19b27(a19b27, a[19], b[27]);
	and and_a19b28(a19b28, a[19], b[28]);
	and and_a19b29(a19b29, a[19], b[29]);
	and and_a19b30(a19b30, a[19], b[30]);
	nand nand_a19b31(not_a19b31, a[19], b[31]);
	and and_a20b0(a20b0, a[20], b[0]);
	and and_a20b1(a20b1, a[20], b[1]);
	and and_a20b2(a20b2, a[20], b[2]);
	and and_a20b3(a20b3, a[20], b[3]);
	and and_a20b4(a20b4, a[20], b[4]);
	and and_a20b5(a20b5, a[20], b[5]);
	and and_a20b6(a20b6, a[20], b[6]);
	and and_a20b7(a20b7, a[20], b[7]);
	and and_a20b8(a20b8, a[20], b[8]);
	and and_a20b9(a20b9, a[20], b[9]);
	and and_a20b10(a20b10, a[20], b[10]);
	and and_a20b11(a20b11, a[20], b[11]);
	and and_a20b12(a20b12, a[20], b[12]);
	and and_a20b13(a20b13, a[20], b[13]);
	and and_a20b14(a20b14, a[20], b[14]);
	and and_a20b15(a20b15, a[20], b[15]);
	and and_a20b16(a20b16, a[20], b[16]);
	and and_a20b17(a20b17, a[20], b[17]);
	and and_a20b18(a20b18, a[20], b[18]);
	and and_a20b19(a20b19, a[20], b[19]);
	and and_a20b20(a20b20, a[20], b[20]);
	and and_a20b21(a20b21, a[20], b[21]);
	and and_a20b22(a20b22, a[20], b[22]);
	and and_a20b23(a20b23, a[20], b[23]);
	and and_a20b24(a20b24, a[20], b[24]);
	and and_a20b25(a20b25, a[20], b[25]);
	and and_a20b26(a20b26, a[20], b[26]);
	and and_a20b27(a20b27, a[20], b[27]);
	and and_a20b28(a20b28, a[20], b[28]);
	and and_a20b29(a20b29, a[20], b[29]);
	and and_a20b30(a20b30, a[20], b[30]);
	nand nand_a20b31(not_a20b31, a[20], b[31]);
	and and_a21b0(a21b0, a[21], b[0]);
	and and_a21b1(a21b1, a[21], b[1]);
	and and_a21b2(a21b2, a[21], b[2]);
	and and_a21b3(a21b3, a[21], b[3]);
	and and_a21b4(a21b4, a[21], b[4]);
	and and_a21b5(a21b5, a[21], b[5]);
	and and_a21b6(a21b6, a[21], b[6]);
	and and_a21b7(a21b7, a[21], b[7]);
	and and_a21b8(a21b8, a[21], b[8]);
	and and_a21b9(a21b9, a[21], b[9]);
	and and_a21b10(a21b10, a[21], b[10]);
	and and_a21b11(a21b11, a[21], b[11]);
	and and_a21b12(a21b12, a[21], b[12]);
	and and_a21b13(a21b13, a[21], b[13]);
	and and_a21b14(a21b14, a[21], b[14]);
	and and_a21b15(a21b15, a[21], b[15]);
	and and_a21b16(a21b16, a[21], b[16]);
	and and_a21b17(a21b17, a[21], b[17]);
	and and_a21b18(a21b18, a[21], b[18]);
	and and_a21b19(a21b19, a[21], b[19]);
	and and_a21b20(a21b20, a[21], b[20]);
	and and_a21b21(a21b21, a[21], b[21]);
	and and_a21b22(a21b22, a[21], b[22]);
	and and_a21b23(a21b23, a[21], b[23]);
	and and_a21b24(a21b24, a[21], b[24]);
	and and_a21b25(a21b25, a[21], b[25]);
	and and_a21b26(a21b26, a[21], b[26]);
	and and_a21b27(a21b27, a[21], b[27]);
	and and_a21b28(a21b28, a[21], b[28]);
	and and_a21b29(a21b29, a[21], b[29]);
	and and_a21b30(a21b30, a[21], b[30]);
	nand nand_a21b31(not_a21b31, a[21], b[31]);
	and and_a22b0(a22b0, a[22], b[0]);
	and and_a22b1(a22b1, a[22], b[1]);
	and and_a22b2(a22b2, a[22], b[2]);
	and and_a22b3(a22b3, a[22], b[3]);
	and and_a22b4(a22b4, a[22], b[4]);
	and and_a22b5(a22b5, a[22], b[5]);
	and and_a22b6(a22b6, a[22], b[6]);
	and and_a22b7(a22b7, a[22], b[7]);
	and and_a22b8(a22b8, a[22], b[8]);
	and and_a22b9(a22b9, a[22], b[9]);
	and and_a22b10(a22b10, a[22], b[10]);
	and and_a22b11(a22b11, a[22], b[11]);
	and and_a22b12(a22b12, a[22], b[12]);
	and and_a22b13(a22b13, a[22], b[13]);
	and and_a22b14(a22b14, a[22], b[14]);
	and and_a22b15(a22b15, a[22], b[15]);
	and and_a22b16(a22b16, a[22], b[16]);
	and and_a22b17(a22b17, a[22], b[17]);
	and and_a22b18(a22b18, a[22], b[18]);
	and and_a22b19(a22b19, a[22], b[19]);
	and and_a22b20(a22b20, a[22], b[20]);
	and and_a22b21(a22b21, a[22], b[21]);
	and and_a22b22(a22b22, a[22], b[22]);
	and and_a22b23(a22b23, a[22], b[23]);
	and and_a22b24(a22b24, a[22], b[24]);
	and and_a22b25(a22b25, a[22], b[25]);
	and and_a22b26(a22b26, a[22], b[26]);
	and and_a22b27(a22b27, a[22], b[27]);
	and and_a22b28(a22b28, a[22], b[28]);
	and and_a22b29(a22b29, a[22], b[29]);
	and and_a22b30(a22b30, a[22], b[30]);
	nand nand_a22b31(not_a22b31, a[22], b[31]);
	and and_a23b0(a23b0, a[23], b[0]);
	and and_a23b1(a23b1, a[23], b[1]);
	and and_a23b2(a23b2, a[23], b[2]);
	and and_a23b3(a23b3, a[23], b[3]);
	and and_a23b4(a23b4, a[23], b[4]);
	and and_a23b5(a23b5, a[23], b[5]);
	and and_a23b6(a23b6, a[23], b[6]);
	and and_a23b7(a23b7, a[23], b[7]);
	and and_a23b8(a23b8, a[23], b[8]);
	and and_a23b9(a23b9, a[23], b[9]);
	and and_a23b10(a23b10, a[23], b[10]);
	and and_a23b11(a23b11, a[23], b[11]);
	and and_a23b12(a23b12, a[23], b[12]);
	and and_a23b13(a23b13, a[23], b[13]);
	and and_a23b14(a23b14, a[23], b[14]);
	and and_a23b15(a23b15, a[23], b[15]);
	and and_a23b16(a23b16, a[23], b[16]);
	and and_a23b17(a23b17, a[23], b[17]);
	and and_a23b18(a23b18, a[23], b[18]);
	and and_a23b19(a23b19, a[23], b[19]);
	and and_a23b20(a23b20, a[23], b[20]);
	and and_a23b21(a23b21, a[23], b[21]);
	and and_a23b22(a23b22, a[23], b[22]);
	and and_a23b23(a23b23, a[23], b[23]);
	and and_a23b24(a23b24, a[23], b[24]);
	and and_a23b25(a23b25, a[23], b[25]);
	and and_a23b26(a23b26, a[23], b[26]);
	and and_a23b27(a23b27, a[23], b[27]);
	and and_a23b28(a23b28, a[23], b[28]);
	and and_a23b29(a23b29, a[23], b[29]);
	and and_a23b30(a23b30, a[23], b[30]);
	nand nand_a23b31(not_a23b31, a[23], b[31]);
	and and_a24b0(a24b0, a[24], b[0]);
	and and_a24b1(a24b1, a[24], b[1]);
	and and_a24b2(a24b2, a[24], b[2]);
	and and_a24b3(a24b3, a[24], b[3]);
	and and_a24b4(a24b4, a[24], b[4]);
	and and_a24b5(a24b5, a[24], b[5]);
	and and_a24b6(a24b6, a[24], b[6]);
	and and_a24b7(a24b7, a[24], b[7]);
	and and_a24b8(a24b8, a[24], b[8]);
	and and_a24b9(a24b9, a[24], b[9]);
	and and_a24b10(a24b10, a[24], b[10]);
	and and_a24b11(a24b11, a[24], b[11]);
	and and_a24b12(a24b12, a[24], b[12]);
	and and_a24b13(a24b13, a[24], b[13]);
	and and_a24b14(a24b14, a[24], b[14]);
	and and_a24b15(a24b15, a[24], b[15]);
	and and_a24b16(a24b16, a[24], b[16]);
	and and_a24b17(a24b17, a[24], b[17]);
	and and_a24b18(a24b18, a[24], b[18]);
	and and_a24b19(a24b19, a[24], b[19]);
	and and_a24b20(a24b20, a[24], b[20]);
	and and_a24b21(a24b21, a[24], b[21]);
	and and_a24b22(a24b22, a[24], b[22]);
	and and_a24b23(a24b23, a[24], b[23]);
	and and_a24b24(a24b24, a[24], b[24]);
	and and_a24b25(a24b25, a[24], b[25]);
	and and_a24b26(a24b26, a[24], b[26]);
	and and_a24b27(a24b27, a[24], b[27]);
	and and_a24b28(a24b28, a[24], b[28]);
	and and_a24b29(a24b29, a[24], b[29]);
	and and_a24b30(a24b30, a[24], b[30]);
	nand nand_a24b31(not_a24b31, a[24], b[31]);
	and and_a25b0(a25b0, a[25], b[0]);
	and and_a25b1(a25b1, a[25], b[1]);
	and and_a25b2(a25b2, a[25], b[2]);
	and and_a25b3(a25b3, a[25], b[3]);
	and and_a25b4(a25b4, a[25], b[4]);
	and and_a25b5(a25b5, a[25], b[5]);
	and and_a25b6(a25b6, a[25], b[6]);
	and and_a25b7(a25b7, a[25], b[7]);
	and and_a25b8(a25b8, a[25], b[8]);
	and and_a25b9(a25b9, a[25], b[9]);
	and and_a25b10(a25b10, a[25], b[10]);
	and and_a25b11(a25b11, a[25], b[11]);
	and and_a25b12(a25b12, a[25], b[12]);
	and and_a25b13(a25b13, a[25], b[13]);
	and and_a25b14(a25b14, a[25], b[14]);
	and and_a25b15(a25b15, a[25], b[15]);
	and and_a25b16(a25b16, a[25], b[16]);
	and and_a25b17(a25b17, a[25], b[17]);
	and and_a25b18(a25b18, a[25], b[18]);
	and and_a25b19(a25b19, a[25], b[19]);
	and and_a25b20(a25b20, a[25], b[20]);
	and and_a25b21(a25b21, a[25], b[21]);
	and and_a25b22(a25b22, a[25], b[22]);
	and and_a25b23(a25b23, a[25], b[23]);
	and and_a25b24(a25b24, a[25], b[24]);
	and and_a25b25(a25b25, a[25], b[25]);
	and and_a25b26(a25b26, a[25], b[26]);
	and and_a25b27(a25b27, a[25], b[27]);
	and and_a25b28(a25b28, a[25], b[28]);
	and and_a25b29(a25b29, a[25], b[29]);
	and and_a25b30(a25b30, a[25], b[30]);
	nand nand_a25b31(not_a25b31, a[25], b[31]);
	and and_a26b0(a26b0, a[26], b[0]);
	and and_a26b1(a26b1, a[26], b[1]);
	and and_a26b2(a26b2, a[26], b[2]);
	and and_a26b3(a26b3, a[26], b[3]);
	and and_a26b4(a26b4, a[26], b[4]);
	and and_a26b5(a26b5, a[26], b[5]);
	and and_a26b6(a26b6, a[26], b[6]);
	and and_a26b7(a26b7, a[26], b[7]);
	and and_a26b8(a26b8, a[26], b[8]);
	and and_a26b9(a26b9, a[26], b[9]);
	and and_a26b10(a26b10, a[26], b[10]);
	and and_a26b11(a26b11, a[26], b[11]);
	and and_a26b12(a26b12, a[26], b[12]);
	and and_a26b13(a26b13, a[26], b[13]);
	and and_a26b14(a26b14, a[26], b[14]);
	and and_a26b15(a26b15, a[26], b[15]);
	and and_a26b16(a26b16, a[26], b[16]);
	and and_a26b17(a26b17, a[26], b[17]);
	and and_a26b18(a26b18, a[26], b[18]);
	and and_a26b19(a26b19, a[26], b[19]);
	and and_a26b20(a26b20, a[26], b[20]);
	and and_a26b21(a26b21, a[26], b[21]);
	and and_a26b22(a26b22, a[26], b[22]);
	and and_a26b23(a26b23, a[26], b[23]);
	and and_a26b24(a26b24, a[26], b[24]);
	and and_a26b25(a26b25, a[26], b[25]);
	and and_a26b26(a26b26, a[26], b[26]);
	and and_a26b27(a26b27, a[26], b[27]);
	and and_a26b28(a26b28, a[26], b[28]);
	and and_a26b29(a26b29, a[26], b[29]);
	and and_a26b30(a26b30, a[26], b[30]);
	nand nand_a26b31(not_a26b31, a[26], b[31]);
	and and_a27b0(a27b0, a[27], b[0]);
	and and_a27b1(a27b1, a[27], b[1]);
	and and_a27b2(a27b2, a[27], b[2]);
	and and_a27b3(a27b3, a[27], b[3]);
	and and_a27b4(a27b4, a[27], b[4]);
	and and_a27b5(a27b5, a[27], b[5]);
	and and_a27b6(a27b6, a[27], b[6]);
	and and_a27b7(a27b7, a[27], b[7]);
	and and_a27b8(a27b8, a[27], b[8]);
	and and_a27b9(a27b9, a[27], b[9]);
	and and_a27b10(a27b10, a[27], b[10]);
	and and_a27b11(a27b11, a[27], b[11]);
	and and_a27b12(a27b12, a[27], b[12]);
	and and_a27b13(a27b13, a[27], b[13]);
	and and_a27b14(a27b14, a[27], b[14]);
	and and_a27b15(a27b15, a[27], b[15]);
	and and_a27b16(a27b16, a[27], b[16]);
	and and_a27b17(a27b17, a[27], b[17]);
	and and_a27b18(a27b18, a[27], b[18]);
	and and_a27b19(a27b19, a[27], b[19]);
	and and_a27b20(a27b20, a[27], b[20]);
	and and_a27b21(a27b21, a[27], b[21]);
	and and_a27b22(a27b22, a[27], b[22]);
	and and_a27b23(a27b23, a[27], b[23]);
	and and_a27b24(a27b24, a[27], b[24]);
	and and_a27b25(a27b25, a[27], b[25]);
	and and_a27b26(a27b26, a[27], b[26]);
	and and_a27b27(a27b27, a[27], b[27]);
	and and_a27b28(a27b28, a[27], b[28]);
	and and_a27b29(a27b29, a[27], b[29]);
	and and_a27b30(a27b30, a[27], b[30]);
	nand nand_a27b31(not_a27b31, a[27], b[31]);
	and and_a28b0(a28b0, a[28], b[0]);
	and and_a28b1(a28b1, a[28], b[1]);
	and and_a28b2(a28b2, a[28], b[2]);
	and and_a28b3(a28b3, a[28], b[3]);
	and and_a28b4(a28b4, a[28], b[4]);
	and and_a28b5(a28b5, a[28], b[5]);
	and and_a28b6(a28b6, a[28], b[6]);
	and and_a28b7(a28b7, a[28], b[7]);
	and and_a28b8(a28b8, a[28], b[8]);
	and and_a28b9(a28b9, a[28], b[9]);
	and and_a28b10(a28b10, a[28], b[10]);
	and and_a28b11(a28b11, a[28], b[11]);
	and and_a28b12(a28b12, a[28], b[12]);
	and and_a28b13(a28b13, a[28], b[13]);
	and and_a28b14(a28b14, a[28], b[14]);
	and and_a28b15(a28b15, a[28], b[15]);
	and and_a28b16(a28b16, a[28], b[16]);
	and and_a28b17(a28b17, a[28], b[17]);
	and and_a28b18(a28b18, a[28], b[18]);
	and and_a28b19(a28b19, a[28], b[19]);
	and and_a28b20(a28b20, a[28], b[20]);
	and and_a28b21(a28b21, a[28], b[21]);
	and and_a28b22(a28b22, a[28], b[22]);
	and and_a28b23(a28b23, a[28], b[23]);
	and and_a28b24(a28b24, a[28], b[24]);
	and and_a28b25(a28b25, a[28], b[25]);
	and and_a28b26(a28b26, a[28], b[26]);
	and and_a28b27(a28b27, a[28], b[27]);
	and and_a28b28(a28b28, a[28], b[28]);
	and and_a28b29(a28b29, a[28], b[29]);
	and and_a28b30(a28b30, a[28], b[30]);
	nand nand_a28b31(not_a28b31, a[28], b[31]);
	and and_a29b0(a29b0, a[29], b[0]);
	and and_a29b1(a29b1, a[29], b[1]);
	and and_a29b2(a29b2, a[29], b[2]);
	and and_a29b3(a29b3, a[29], b[3]);
	and and_a29b4(a29b4, a[29], b[4]);
	and and_a29b5(a29b5, a[29], b[5]);
	and and_a29b6(a29b6, a[29], b[6]);
	and and_a29b7(a29b7, a[29], b[7]);
	and and_a29b8(a29b8, a[29], b[8]);
	and and_a29b9(a29b9, a[29], b[9]);
	and and_a29b10(a29b10, a[29], b[10]);
	and and_a29b11(a29b11, a[29], b[11]);
	and and_a29b12(a29b12, a[29], b[12]);
	and and_a29b13(a29b13, a[29], b[13]);
	and and_a29b14(a29b14, a[29], b[14]);
	and and_a29b15(a29b15, a[29], b[15]);
	and and_a29b16(a29b16, a[29], b[16]);
	and and_a29b17(a29b17, a[29], b[17]);
	and and_a29b18(a29b18, a[29], b[18]);
	and and_a29b19(a29b19, a[29], b[19]);
	and and_a29b20(a29b20, a[29], b[20]);
	and and_a29b21(a29b21, a[29], b[21]);
	and and_a29b22(a29b22, a[29], b[22]);
	and and_a29b23(a29b23, a[29], b[23]);
	and and_a29b24(a29b24, a[29], b[24]);
	and and_a29b25(a29b25, a[29], b[25]);
	and and_a29b26(a29b26, a[29], b[26]);
	and and_a29b27(a29b27, a[29], b[27]);
	and and_a29b28(a29b28, a[29], b[28]);
	and and_a29b29(a29b29, a[29], b[29]);
	and and_a29b30(a29b30, a[29], b[30]);
	nand nand_a29b31(not_a29b31, a[29], b[31]);
	and and_a30b0(a30b0, a[30], b[0]);
	and and_a30b1(a30b1, a[30], b[1]);
	and and_a30b2(a30b2, a[30], b[2]);
	and and_a30b3(a30b3, a[30], b[3]);
	and and_a30b4(a30b4, a[30], b[4]);
	and and_a30b5(a30b5, a[30], b[5]);
	and and_a30b6(a30b6, a[30], b[6]);
	and and_a30b7(a30b7, a[30], b[7]);
	and and_a30b8(a30b8, a[30], b[8]);
	and and_a30b9(a30b9, a[30], b[9]);
	and and_a30b10(a30b10, a[30], b[10]);
	and and_a30b11(a30b11, a[30], b[11]);
	and and_a30b12(a30b12, a[30], b[12]);
	and and_a30b13(a30b13, a[30], b[13]);
	and and_a30b14(a30b14, a[30], b[14]);
	and and_a30b15(a30b15, a[30], b[15]);
	and and_a30b16(a30b16, a[30], b[16]);
	and and_a30b17(a30b17, a[30], b[17]);
	and and_a30b18(a30b18, a[30], b[18]);
	and and_a30b19(a30b19, a[30], b[19]);
	and and_a30b20(a30b20, a[30], b[20]);
	and and_a30b21(a30b21, a[30], b[21]);
	and and_a30b22(a30b22, a[30], b[22]);
	and and_a30b23(a30b23, a[30], b[23]);
	and and_a30b24(a30b24, a[30], b[24]);
	and and_a30b25(a30b25, a[30], b[25]);
	and and_a30b26(a30b26, a[30], b[26]);
	and and_a30b27(a30b27, a[30], b[27]);
	and and_a30b28(a30b28, a[30], b[28]);
	and and_a30b29(a30b29, a[30], b[29]);
	and and_a30b30(a30b30, a[30], b[30]);
	nand nand_a30b31(not_a30b31, a[30], b[31]);
	nand nand_a31b0(not_a31b0, a[31], b[0]);
	nand nand_a31b1(not_a31b1, a[31], b[1]);
	nand nand_a31b2(not_a31b2, a[31], b[2]);
	nand nand_a31b3(not_a31b3, a[31], b[3]);
	nand nand_a31b4(not_a31b4, a[31], b[4]);
	nand nand_a31b5(not_a31b5, a[31], b[5]);
	nand nand_a31b6(not_a31b6, a[31], b[6]);
	nand nand_a31b7(not_a31b7, a[31], b[7]);
	nand nand_a31b8(not_a31b8, a[31], b[8]);
	nand nand_a31b9(not_a31b9, a[31], b[9]);
	nand nand_a31b10(not_a31b10, a[31], b[10]);
	nand nand_a31b11(not_a31b11, a[31], b[11]);
	nand nand_a31b12(not_a31b12, a[31], b[12]);
	nand nand_a31b13(not_a31b13, a[31], b[13]);
	nand nand_a31b14(not_a31b14, a[31], b[14]);
	nand nand_a31b15(not_a31b15, a[31], b[15]);
	nand nand_a31b16(not_a31b16, a[31], b[16]);
	nand nand_a31b17(not_a31b17, a[31], b[17]);
	nand nand_a31b18(not_a31b18, a[31], b[18]);
	nand nand_a31b19(not_a31b19, a[31], b[19]);
	nand nand_a31b20(not_a31b20, a[31], b[20]);
	nand nand_a31b21(not_a31b21, a[31], b[21]);
	nand nand_a31b22(not_a31b22, a[31], b[22]);
	nand nand_a31b23(not_a31b23, a[31], b[23]);
	nand nand_a31b24(not_a31b24, a[31], b[24]);
	nand nand_a31b25(not_a31b25, a[31], b[25]);
	nand nand_a31b26(not_a31b26, a[31], b[26]);
	nand nand_a31b27(not_a31b27, a[31], b[27]);
	nand nand_a31b28(not_a31b28, a[31], b[28]);
	nand nand_a31b29(not_a31b29, a[31], b[29]);
	nand nand_a31b30(not_a31b30, a[31], b[30]);
	and and_a31b31(a31b31, a[31], b[31]);
	half_adder (a0b1, a1b0, w_1_1_1, w_1_2_1);
	full_adder (a0b2, a1b1, a2b0, w_1_2_2, w_1_3_1);
	full_adder (a0b3, a1b2, a2b1, w_1_3_2, w_1_4_1);
	full_adder (a0b4, a1b3, a2b2, w_1_4_2, w_1_5_1);
	half_adder (a3b1, a4b0, w_1_4_3, w_1_5_2);
	full_adder (a0b5, a1b4, a2b3, w_1_5_3, w_1_6_1);
	full_adder (a3b2, a4b1, a5b0, w_1_5_4, w_1_6_2);
	full_adder (a0b6, a1b5, a2b4, w_1_6_3, w_1_7_1);
	full_adder (a3b3, a4b2, a5b1, w_1_6_4, w_1_7_2);
	full_adder (a0b7, a1b6, a2b5, w_1_7_3, w_1_8_1);
	full_adder (a3b4, a4b3, a5b2, w_1_7_4, w_1_8_2);
	half_adder (a6b1, a7b0, w_1_7_5, w_1_8_3);
	full_adder (a0b8, a1b7, a2b6, w_1_8_4, w_1_9_1);
	full_adder (a3b5, a4b4, a5b3, w_1_8_5, w_1_9_2);
	full_adder (a6b2, a7b1, a8b0, w_1_8_6, w_1_9_3);
	full_adder (a0b9, a1b8, a2b7, w_1_9_4, w_1_10_1);
	full_adder (a3b6, a4b5, a5b4, w_1_9_5, w_1_10_2);
	full_adder (a6b3, a7b2, a8b1, w_1_9_6, w_1_10_3);
	full_adder (a0b10, a1b9, a2b8, w_1_10_4, w_1_11_1);
	full_adder (a3b7, a4b6, a5b5, w_1_10_5, w_1_11_2);
	full_adder (a6b4, a7b3, a8b2, w_1_10_6, w_1_11_3);
	half_adder (a9b1, a10b0, w_1_10_7, w_1_11_4);
	full_adder (a0b11, a1b10, a2b9, w_1_11_5, w_1_12_1);
	full_adder (a3b8, a4b7, a5b6, w_1_11_6, w_1_12_2);
	full_adder (a6b5, a7b4, a8b3, w_1_11_7, w_1_12_3);
	full_adder (a9b2, a10b1, a11b0, w_1_11_8, w_1_12_4);
	full_adder (a0b12, a1b11, a2b10, w_1_12_5, w_1_13_1);
	full_adder (a3b9, a4b8, a5b7, w_1_12_6, w_1_13_2);
	full_adder (a6b6, a7b5, a8b4, w_1_12_7, w_1_13_3);
	full_adder (a9b3, a10b2, a11b1, w_1_12_8, w_1_13_4);
	full_adder (a0b13, a1b12, a2b11, w_1_13_5, w_1_14_1);
	full_adder (a3b10, a4b9, a5b8, w_1_13_6, w_1_14_2);
	full_adder (a6b7, a7b6, a8b5, w_1_13_7, w_1_14_3);
	full_adder (a9b4, a10b3, a11b2, w_1_13_8, w_1_14_4);
	half_adder (a12b1, a13b0, w_1_13_9, w_1_14_5);
	full_adder (a0b14, a1b13, a2b12, w_1_14_6, w_1_15_1);
	full_adder (a3b11, a4b10, a5b9, w_1_14_7, w_1_15_2);
	full_adder (a6b8, a7b7, a8b6, w_1_14_8, w_1_15_3);
	full_adder (a9b5, a10b4, a11b3, w_1_14_9, w_1_15_4);
	full_adder (a12b2, a13b1, a14b0, w_1_14_10, w_1_15_5);
	full_adder (a0b15, a1b14, a2b13, w_1_15_6, w_1_16_1);
	full_adder (a3b12, a4b11, a5b10, w_1_15_7, w_1_16_2);
	full_adder (a6b9, a7b8, a8b7, w_1_15_8, w_1_16_3);
	full_adder (a9b6, a10b5, a11b4, w_1_15_9, w_1_16_4);
	full_adder (a12b3, a13b2, a14b1, w_1_15_10, w_1_16_5);
	full_adder (a0b16, a1b15, a2b14, w_1_16_6, w_1_17_1);
	full_adder (a3b13, a4b12, a5b11, w_1_16_7, w_1_17_2);
	full_adder (a6b10, a7b9, a8b8, w_1_16_8, w_1_17_3);
	full_adder (a9b7, a10b6, a11b5, w_1_16_9, w_1_17_4);
	full_adder (a12b4, a13b3, a14b2, w_1_16_10, w_1_17_5);
	half_adder (a15b1, a16b0, w_1_16_11, w_1_17_6);
	full_adder (a0b17, a1b16, a2b15, w_1_17_7, w_1_18_1);
	full_adder (a3b14, a4b13, a5b12, w_1_17_8, w_1_18_2);
	full_adder (a6b11, a7b10, a8b9, w_1_17_9, w_1_18_3);
	full_adder (a9b8, a10b7, a11b6, w_1_17_10, w_1_18_4);
	full_adder (a12b5, a13b4, a14b3, w_1_17_11, w_1_18_5);
	full_adder (a15b2, a16b1, a17b0, w_1_17_12, w_1_18_6);
	full_adder (a0b18, a1b17, a2b16, w_1_18_7, w_1_19_1);
	full_adder (a3b15, a4b14, a5b13, w_1_18_8, w_1_19_2);
	full_adder (a6b12, a7b11, a8b10, w_1_18_9, w_1_19_3);
	full_adder (a9b9, a10b8, a11b7, w_1_18_10, w_1_19_4);
	full_adder (a12b6, a13b5, a14b4, w_1_18_11, w_1_19_5);
	full_adder (a15b3, a16b2, a17b1, w_1_18_12, w_1_19_6);
	full_adder (a0b19, a1b18, a2b17, w_1_19_7, w_1_20_1);
	full_adder (a3b16, a4b15, a5b14, w_1_19_8, w_1_20_2);
	full_adder (a6b13, a7b12, a8b11, w_1_19_9, w_1_20_3);
	full_adder (a9b10, a10b9, a11b8, w_1_19_10, w_1_20_4);
	full_adder (a12b7, a13b6, a14b5, w_1_19_11, w_1_20_5);
	full_adder (a15b4, a16b3, a17b2, w_1_19_12, w_1_20_6);
	half_adder (a18b1, a19b0, w_1_19_13, w_1_20_7);
	full_adder (a0b20, a1b19, a2b18, w_1_20_8, w_1_21_1);
	full_adder (a3b17, a4b16, a5b15, w_1_20_9, w_1_21_2);
	full_adder (a6b14, a7b13, a8b12, w_1_20_10, w_1_21_3);
	full_adder (a9b11, a10b10, a11b9, w_1_20_11, w_1_21_4);
	full_adder (a12b8, a13b7, a14b6, w_1_20_12, w_1_21_5);
	full_adder (a15b5, a16b4, a17b3, w_1_20_13, w_1_21_6);
	full_adder (a18b2, a19b1, a20b0, w_1_20_14, w_1_21_7);
	full_adder (a0b21, a1b20, a2b19, w_1_21_8, w_1_22_1);
	full_adder (a3b18, a4b17, a5b16, w_1_21_9, w_1_22_2);
	full_adder (a6b15, a7b14, a8b13, w_1_21_10, w_1_22_3);
	full_adder (a9b12, a10b11, a11b10, w_1_21_11, w_1_22_4);
	full_adder (a12b9, a13b8, a14b7, w_1_21_12, w_1_22_5);
	full_adder (a15b6, a16b5, a17b4, w_1_21_13, w_1_22_6);
	full_adder (a18b3, a19b2, a20b1, w_1_21_14, w_1_22_7);
	full_adder (a0b22, a1b21, a2b20, w_1_22_8, w_1_23_1);
	full_adder (a3b19, a4b18, a5b17, w_1_22_9, w_1_23_2);
	full_adder (a6b16, a7b15, a8b14, w_1_22_10, w_1_23_3);
	full_adder (a9b13, a10b12, a11b11, w_1_22_11, w_1_23_4);
	full_adder (a12b10, a13b9, a14b8, w_1_22_12, w_1_23_5);
	full_adder (a15b7, a16b6, a17b5, w_1_22_13, w_1_23_6);
	full_adder (a18b4, a19b3, a20b2, w_1_22_14, w_1_23_7);
	half_adder (a21b1, a22b0, w_1_22_15, w_1_23_8);
	full_adder (a0b23, a1b22, a2b21, w_1_23_9, w_1_24_1);
	full_adder (a3b20, a4b19, a5b18, w_1_23_10, w_1_24_2);
	full_adder (a6b17, a7b16, a8b15, w_1_23_11, w_1_24_3);
	full_adder (a9b14, a10b13, a11b12, w_1_23_12, w_1_24_4);
	full_adder (a12b11, a13b10, a14b9, w_1_23_13, w_1_24_5);
	full_adder (a15b8, a16b7, a17b6, w_1_23_14, w_1_24_6);
	full_adder (a18b5, a19b4, a20b3, w_1_23_15, w_1_24_7);
	full_adder (a21b2, a22b1, a23b0, w_1_23_16, w_1_24_8);
	full_adder (a0b24, a1b23, a2b22, w_1_24_9, w_1_25_1);
	full_adder (a3b21, a4b20, a5b19, w_1_24_10, w_1_25_2);
	full_adder (a6b18, a7b17, a8b16, w_1_24_11, w_1_25_3);
	full_adder (a9b15, a10b14, a11b13, w_1_24_12, w_1_25_4);
	full_adder (a12b12, a13b11, a14b10, w_1_24_13, w_1_25_5);
	full_adder (a15b9, a16b8, a17b7, w_1_24_14, w_1_25_6);
	full_adder (a18b6, a19b5, a20b4, w_1_24_15, w_1_25_7);
	full_adder (a21b3, a22b2, a23b1, w_1_24_16, w_1_25_8);
	full_adder (a0b25, a1b24, a2b23, w_1_25_9, w_1_26_1);
	full_adder (a3b22, a4b21, a5b20, w_1_25_10, w_1_26_2);
	full_adder (a6b19, a7b18, a8b17, w_1_25_11, w_1_26_3);
	full_adder (a9b16, a10b15, a11b14, w_1_25_12, w_1_26_4);
	full_adder (a12b13, a13b12, a14b11, w_1_25_13, w_1_26_5);
	full_adder (a15b10, a16b9, a17b8, w_1_25_14, w_1_26_6);
	full_adder (a18b7, a19b6, a20b5, w_1_25_15, w_1_26_7);
	full_adder (a21b4, a22b3, a23b2, w_1_25_16, w_1_26_8);
	half_adder (a24b1, a25b0, w_1_25_17, w_1_26_9);
	full_adder (a0b26, a1b25, a2b24, w_1_26_10, w_1_27_1);
	full_adder (a3b23, a4b22, a5b21, w_1_26_11, w_1_27_2);
	full_adder (a6b20, a7b19, a8b18, w_1_26_12, w_1_27_3);
	full_adder (a9b17, a10b16, a11b15, w_1_26_13, w_1_27_4);
	full_adder (a12b14, a13b13, a14b12, w_1_26_14, w_1_27_5);
	full_adder (a15b11, a16b10, a17b9, w_1_26_15, w_1_27_6);
	full_adder (a18b8, a19b7, a20b6, w_1_26_16, w_1_27_7);
	full_adder (a21b5, a22b4, a23b3, w_1_26_17, w_1_27_8);
	full_adder (a24b2, a25b1, a26b0, w_1_26_18, w_1_27_9);
	full_adder (a0b27, a1b26, a2b25, w_1_27_10, w_1_28_1);
	full_adder (a3b24, a4b23, a5b22, w_1_27_11, w_1_28_2);
	full_adder (a6b21, a7b20, a8b19, w_1_27_12, w_1_28_3);
	full_adder (a9b18, a10b17, a11b16, w_1_27_13, w_1_28_4);
	full_adder (a12b15, a13b14, a14b13, w_1_27_14, w_1_28_5);
	full_adder (a15b12, a16b11, a17b10, w_1_27_15, w_1_28_6);
	full_adder (a18b9, a19b8, a20b7, w_1_27_16, w_1_28_7);
	full_adder (a21b6, a22b5, a23b4, w_1_27_17, w_1_28_8);
	full_adder (a24b3, a25b2, a26b1, w_1_27_18, w_1_28_9);
	full_adder (a0b28, a1b27, a2b26, w_1_28_10, w_1_29_1);
	full_adder (a3b25, a4b24, a5b23, w_1_28_11, w_1_29_2);
	full_adder (a6b22, a7b21, a8b20, w_1_28_12, w_1_29_3);
	full_adder (a9b19, a10b18, a11b17, w_1_28_13, w_1_29_4);
	full_adder (a12b16, a13b15, a14b14, w_1_28_14, w_1_29_5);
	full_adder (a15b13, a16b12, a17b11, w_1_28_15, w_1_29_6);
	full_adder (a18b10, a19b9, a20b8, w_1_28_16, w_1_29_7);
	full_adder (a21b7, a22b6, a23b5, w_1_28_17, w_1_29_8);
	full_adder (a24b4, a25b3, a26b2, w_1_28_18, w_1_29_9);
	half_adder (a27b1, a28b0, w_1_28_19, w_1_29_10);
	full_adder (a0b29, a1b28, a2b27, w_1_29_11, w_1_30_1);
	full_adder (a3b26, a4b25, a5b24, w_1_29_12, w_1_30_2);
	full_adder (a6b23, a7b22, a8b21, w_1_29_13, w_1_30_3);
	full_adder (a9b20, a10b19, a11b18, w_1_29_14, w_1_30_4);
	full_adder (a12b17, a13b16, a14b15, w_1_29_15, w_1_30_5);
	full_adder (a15b14, a16b13, a17b12, w_1_29_16, w_1_30_6);
	full_adder (a18b11, a19b10, a20b9, w_1_29_17, w_1_30_7);
	full_adder (a21b8, a22b7, a23b6, w_1_29_18, w_1_30_8);
	full_adder (a24b5, a25b4, a26b3, w_1_29_19, w_1_30_9);
	full_adder (a27b2, a28b1, a29b0, w_1_29_20, w_1_30_10);
	full_adder (a0b30, a1b29, a2b28, w_1_30_11, w_1_31_1);
	full_adder (a3b27, a4b26, a5b25, w_1_30_12, w_1_31_2);
	full_adder (a6b24, a7b23, a8b22, w_1_30_13, w_1_31_3);
	full_adder (a9b21, a10b20, a11b19, w_1_30_14, w_1_31_4);
	full_adder (a12b18, a13b17, a14b16, w_1_30_15, w_1_31_5);
	full_adder (a15b15, a16b14, a17b13, w_1_30_16, w_1_31_6);
	full_adder (a18b12, a19b11, a20b10, w_1_30_17, w_1_31_7);
	full_adder (a21b9, a22b8, a23b7, w_1_30_18, w_1_31_8);
	full_adder (a24b6, a25b5, a26b4, w_1_30_19, w_1_31_9);
	full_adder (a27b3, a28b2, a29b1, w_1_30_20, w_1_31_10);
	full_adder (not_a0b31, a1b30, a2b29, w_1_31_11, w_1_32_1);
	full_adder (a3b28, a4b27, a5b26, w_1_31_12, w_1_32_2);
	full_adder (a6b25, a7b24, a8b23, w_1_31_13, w_1_32_3);
	full_adder (a9b22, a10b21, a11b20, w_1_31_14, w_1_32_4);
	full_adder (a12b19, a13b18, a14b17, w_1_31_15, w_1_32_5);
	full_adder (a15b16, a16b15, a17b14, w_1_31_16, w_1_32_6);
	full_adder (a18b13, a19b12, a20b11, w_1_31_17, w_1_32_7);
	full_adder (a21b10, a22b9, a23b8, w_1_31_18, w_1_32_8);
	full_adder (a24b7, a25b6, a26b5, w_1_31_19, w_1_32_9);
	full_adder (a27b4, a28b3, a29b2, w_1_31_20, w_1_32_10);
	half_adder (a30b1, not_a31b0, w_1_31_21, w_1_32_11);
	full_adder (not_a1b31, a2b30, a3b29, w_1_32_12, w_1_33_1);
	full_adder (a4b28, a5b27, a6b26, w_1_32_13, w_1_33_2);
	full_adder (a7b25, a8b24, a9b23, w_1_32_14, w_1_33_3);
	full_adder (a10b22, a11b21, a12b20, w_1_32_15, w_1_33_4);
	full_adder (a13b19, a14b18, a15b17, w_1_32_16, w_1_33_5);
	full_adder (a16b16, a17b15, a18b14, w_1_32_17, w_1_33_6);
	full_adder (a19b13, a20b12, a21b11, w_1_32_18, w_1_33_7);
	full_adder (a22b10, a23b9, a24b8, w_1_32_19, w_1_33_8);
	full_adder (a25b7, a26b6, a27b5, w_1_32_20, w_1_33_9);
	full_adder (a28b4, a29b3, a30b2, w_1_32_21, w_1_33_10);
	half_adder (not_a31b1, 1, w_1_32_22, w_1_33_11);
	full_adder (not_a2b31, a3b30, a4b29, w_1_33_12, w_1_34_1);
	full_adder (a5b28, a6b27, a7b26, w_1_33_13, w_1_34_2);
	full_adder (a8b25, a9b24, a10b23, w_1_33_14, w_1_34_3);
	full_adder (a11b22, a12b21, a13b20, w_1_33_15, w_1_34_4);
	full_adder (a14b19, a15b18, a16b17, w_1_33_16, w_1_34_5);
	full_adder (a17b16, a18b15, a19b14, w_1_33_17, w_1_34_6);
	full_adder (a20b13, a21b12, a22b11, w_1_33_18, w_1_34_7);
	full_adder (a23b10, a24b9, a25b8, w_1_33_19, w_1_34_8);
	full_adder (a26b7, a27b6, a28b5, w_1_33_20, w_1_34_9);
	full_adder (a29b4, a30b3, not_a31b2, w_1_33_21, w_1_34_10);
	full_adder (not_a3b31, a4b30, a5b29, w_1_34_11, w_1_35_1);
	full_adder (a6b28, a7b27, a8b26, w_1_34_12, w_1_35_2);
	full_adder (a9b25, a10b24, a11b23, w_1_34_13, w_1_35_3);
	full_adder (a12b22, a13b21, a14b20, w_1_34_14, w_1_35_4);
	full_adder (a15b19, a16b18, a17b17, w_1_34_15, w_1_35_5);
	full_adder (a18b16, a19b15, a20b14, w_1_34_16, w_1_35_6);
	full_adder (a21b13, a22b12, a23b11, w_1_34_17, w_1_35_7);
	full_adder (a24b10, a25b9, a26b8, w_1_34_18, w_1_35_8);
	full_adder (a27b7, a28b6, a29b5, w_1_34_19, w_1_35_9);
	half_adder (a30b4, not_a31b3, w_1_34_20, w_1_35_10);
	full_adder (not_a4b31, a5b30, a6b29, w_1_35_11, w_1_36_1);
	full_adder (a7b28, a8b27, a9b26, w_1_35_12, w_1_36_2);
	full_adder (a10b25, a11b24, a12b23, w_1_35_13, w_1_36_3);
	full_adder (a13b22, a14b21, a15b20, w_1_35_14, w_1_36_4);
	full_adder (a16b19, a17b18, a18b17, w_1_35_15, w_1_36_5);
	full_adder (a19b16, a20b15, a21b14, w_1_35_16, w_1_36_6);
	full_adder (a22b13, a23b12, a24b11, w_1_35_17, w_1_36_7);
	full_adder (a25b10, a26b9, a27b8, w_1_35_18, w_1_36_8);
	full_adder (a28b7, a29b6, a30b5, w_1_35_19, w_1_36_9);
	full_adder (not_a5b31, a6b30, a7b29, w_1_36_10, w_1_37_1);
	full_adder (a8b28, a9b27, a10b26, w_1_36_11, w_1_37_2);
	full_adder (a11b25, a12b24, a13b23, w_1_36_12, w_1_37_3);
	full_adder (a14b22, a15b21, a16b20, w_1_36_13, w_1_37_4);
	full_adder (a17b19, a18b18, a19b17, w_1_36_14, w_1_37_5);
	full_adder (a20b16, a21b15, a22b14, w_1_36_15, w_1_37_6);
	full_adder (a23b13, a24b12, a25b11, w_1_36_16, w_1_37_7);
	full_adder (a26b10, a27b9, a28b8, w_1_36_17, w_1_37_8);
	full_adder (a29b7, a30b6, not_a31b5, w_1_36_18, w_1_37_9);
	full_adder (not_a6b31, a7b30, a8b29, w_1_37_10, w_1_38_1);
	full_adder (a9b28, a10b27, a11b26, w_1_37_11, w_1_38_2);
	full_adder (a12b25, a13b24, a14b23, w_1_37_12, w_1_38_3);
	full_adder (a15b22, a16b21, a17b20, w_1_37_13, w_1_38_4);
	full_adder (a18b19, a19b18, a20b17, w_1_37_14, w_1_38_5);
	full_adder (a21b16, a22b15, a23b14, w_1_37_15, w_1_38_6);
	full_adder (a24b13, a25b12, a26b11, w_1_37_16, w_1_38_7);
	full_adder (a27b10, a28b9, a29b8, w_1_37_17, w_1_38_8);
	half_adder (a30b7, not_a31b6, w_1_37_18, w_1_38_9);
	full_adder (not_a7b31, a8b30, a9b29, w_1_38_10, w_1_39_1);
	full_adder (a10b28, a11b27, a12b26, w_1_38_11, w_1_39_2);
	full_adder (a13b25, a14b24, a15b23, w_1_38_12, w_1_39_3);
	full_adder (a16b22, a17b21, a18b20, w_1_38_13, w_1_39_4);
	full_adder (a19b19, a20b18, a21b17, w_1_38_14, w_1_39_5);
	full_adder (a22b16, a23b15, a24b14, w_1_38_15, w_1_39_6);
	full_adder (a25b13, a26b12, a27b11, w_1_38_16, w_1_39_7);
	full_adder (a28b10, a29b9, a30b8, w_1_38_17, w_1_39_8);
	full_adder (not_a8b31, a9b30, a10b29, w_1_39_9, w_1_40_1);
	full_adder (a11b28, a12b27, a13b26, w_1_39_10, w_1_40_2);
	full_adder (a14b25, a15b24, a16b23, w_1_39_11, w_1_40_3);
	full_adder (a17b22, a18b21, a19b20, w_1_39_12, w_1_40_4);
	full_adder (a20b19, a21b18, a22b17, w_1_39_13, w_1_40_5);
	full_adder (a23b16, a24b15, a25b14, w_1_39_14, w_1_40_6);
	full_adder (a26b13, a27b12, a28b11, w_1_39_15, w_1_40_7);
	full_adder (a29b10, a30b9, not_a31b8, w_1_39_16, w_1_40_8);
	full_adder (not_a9b31, a10b30, a11b29, w_1_40_9, w_1_41_1);
	full_adder (a12b28, a13b27, a14b26, w_1_40_10, w_1_41_2);
	full_adder (a15b25, a16b24, a17b23, w_1_40_11, w_1_41_3);
	full_adder (a18b22, a19b21, a20b20, w_1_40_12, w_1_41_4);
	full_adder (a21b19, a22b18, a23b17, w_1_40_13, w_1_41_5);
	full_adder (a24b16, a25b15, a26b14, w_1_40_14, w_1_41_6);
	full_adder (a27b13, a28b12, a29b11, w_1_40_15, w_1_41_7);
	half_adder (a30b10, not_a31b9, w_1_40_16, w_1_41_8);
	full_adder (not_a10b31, a11b30, a12b29, w_1_41_9, w_1_42_1);
	full_adder (a13b28, a14b27, a15b26, w_1_41_10, w_1_42_2);
	full_adder (a16b25, a17b24, a18b23, w_1_41_11, w_1_42_3);
	full_adder (a19b22, a20b21, a21b20, w_1_41_12, w_1_42_4);
	full_adder (a22b19, a23b18, a24b17, w_1_41_13, w_1_42_5);
	full_adder (a25b16, a26b15, a27b14, w_1_41_14, w_1_42_6);
	full_adder (a28b13, a29b12, a30b11, w_1_41_15, w_1_42_7);
	full_adder (not_a11b31, a12b30, a13b29, w_1_42_8, w_1_43_1);
	full_adder (a14b28, a15b27, a16b26, w_1_42_9, w_1_43_2);
	full_adder (a17b25, a18b24, a19b23, w_1_42_10, w_1_43_3);
	full_adder (a20b22, a21b21, a22b20, w_1_42_11, w_1_43_4);
	full_adder (a23b19, a24b18, a25b17, w_1_42_12, w_1_43_5);
	full_adder (a26b16, a27b15, a28b14, w_1_42_13, w_1_43_6);
	full_adder (a29b13, a30b12, not_a31b11, w_1_42_14, w_1_43_7);
	full_adder (not_a12b31, a13b30, a14b29, w_1_43_8, w_1_44_1);
	full_adder (a15b28, a16b27, a17b26, w_1_43_9, w_1_44_2);
	full_adder (a18b25, a19b24, a20b23, w_1_43_10, w_1_44_3);
	full_adder (a21b22, a22b21, a23b20, w_1_43_11, w_1_44_4);
	full_adder (a24b19, a25b18, a26b17, w_1_43_12, w_1_44_5);
	full_adder (a27b16, a28b15, a29b14, w_1_43_13, w_1_44_6);
	half_adder (a30b13, not_a31b12, w_1_43_14, w_1_44_7);
	full_adder (not_a13b31, a14b30, a15b29, w_1_44_8, w_1_45_1);
	full_adder (a16b28, a17b27, a18b26, w_1_44_9, w_1_45_2);
	full_adder (a19b25, a20b24, a21b23, w_1_44_10, w_1_45_3);
	full_adder (a22b22, a23b21, a24b20, w_1_44_11, w_1_45_4);
	full_adder (a25b19, a26b18, a27b17, w_1_44_12, w_1_45_5);
	full_adder (a28b16, a29b15, a30b14, w_1_44_13, w_1_45_6);
	full_adder (not_a14b31, a15b30, a16b29, w_1_45_7, w_1_46_1);
	full_adder (a17b28, a18b27, a19b26, w_1_45_8, w_1_46_2);
	full_adder (a20b25, a21b24, a22b23, w_1_45_9, w_1_46_3);
	full_adder (a23b22, a24b21, a25b20, w_1_45_10, w_1_46_4);
	full_adder (a26b19, a27b18, a28b17, w_1_45_11, w_1_46_5);
	full_adder (a29b16, a30b15, not_a31b14, w_1_45_12, w_1_46_6);
	full_adder (not_a15b31, a16b30, a17b29, w_1_46_7, w_1_47_1);
	full_adder (a18b28, a19b27, a20b26, w_1_46_8, w_1_47_2);
	full_adder (a21b25, a22b24, a23b23, w_1_46_9, w_1_47_3);
	full_adder (a24b22, a25b21, a26b20, w_1_46_10, w_1_47_4);
	full_adder (a27b19, a28b18, a29b17, w_1_46_11, w_1_47_5);
	half_adder (a30b16, not_a31b15, w_1_46_12, w_1_47_6);
	full_adder (not_a16b31, a17b30, a18b29, w_1_47_7, w_1_48_1);
	full_adder (a19b28, a20b27, a21b26, w_1_47_8, w_1_48_2);
	full_adder (a22b25, a23b24, a24b23, w_1_47_9, w_1_48_3);
	full_adder (a25b22, a26b21, a27b20, w_1_47_10, w_1_48_4);
	full_adder (a28b19, a29b18, a30b17, w_1_47_11, w_1_48_5);
	full_adder (not_a17b31, a18b30, a19b29, w_1_48_6, w_1_49_1);
	full_adder (a20b28, a21b27, a22b26, w_1_48_7, w_1_49_2);
	full_adder (a23b25, a24b24, a25b23, w_1_48_8, w_1_49_3);
	full_adder (a26b22, a27b21, a28b20, w_1_48_9, w_1_49_4);
	full_adder (a29b19, a30b18, not_a31b17, w_1_48_10, w_1_49_5);
	full_adder (not_a18b31, a19b30, a20b29, w_1_49_6, w_1_50_1);
	full_adder (a21b28, a22b27, a23b26, w_1_49_7, w_1_50_2);
	full_adder (a24b25, a25b24, a26b23, w_1_49_8, w_1_50_3);
	full_adder (a27b22, a28b21, a29b20, w_1_49_9, w_1_50_4);
	half_adder (a30b19, not_a31b18, w_1_49_10, w_1_50_5);
	full_adder (not_a19b31, a20b30, a21b29, w_1_50_6, w_1_51_1);
	full_adder (a22b28, a23b27, a24b26, w_1_50_7, w_1_51_2);
	full_adder (a25b25, a26b24, a27b23, w_1_50_8, w_1_51_3);
	full_adder (a28b22, a29b21, a30b20, w_1_50_9, w_1_51_4);
	full_adder (not_a20b31, a21b30, a22b29, w_1_51_5, w_1_52_1);
	full_adder (a23b28, a24b27, a25b26, w_1_51_6, w_1_52_2);
	full_adder (a26b25, a27b24, a28b23, w_1_51_7, w_1_52_3);
	full_adder (a29b22, a30b21, not_a31b20, w_1_51_8, w_1_52_4);
	full_adder (not_a21b31, a22b30, a23b29, w_1_52_5, w_1_53_1);
	full_adder (a24b28, a25b27, a26b26, w_1_52_6, w_1_53_2);
	full_adder (a27b25, a28b24, a29b23, w_1_52_7, w_1_53_3);
	half_adder (a30b22, not_a31b21, w_1_52_8, w_1_53_4);
	full_adder (not_a22b31, a23b30, a24b29, w_1_53_5, w_1_54_1);
	full_adder (a25b28, a26b27, a27b26, w_1_53_6, w_1_54_2);
	full_adder (a28b25, a29b24, a30b23, w_1_53_7, w_1_54_3);
	full_adder (not_a23b31, a24b30, a25b29, w_1_54_4, w_1_55_1);
	full_adder (a26b28, a27b27, a28b26, w_1_54_5, w_1_55_2);
	full_adder (a29b25, a30b24, not_a31b23, w_1_54_6, w_1_55_3);
	full_adder (not_a24b31, a25b30, a26b29, w_1_55_4, w_1_56_1);
	full_adder (a27b28, a28b27, a29b26, w_1_55_5, w_1_56_2);
	half_adder (a30b25, not_a31b24, w_1_55_6, w_1_56_3);
	full_adder (not_a25b31, a26b30, a27b29, w_1_56_4, w_1_57_1);
	full_adder (a28b28, a29b27, a30b26, w_1_56_5, w_1_57_2);
	full_adder (not_a26b31, a27b30, a28b29, w_1_57_3, w_1_58_1);
	full_adder (a29b28, a30b27, not_a31b26, w_1_57_4, w_1_58_2);
	full_adder (not_a27b31, a28b30, a29b29, w_1_58_3, w_1_59_1);
	half_adder (a30b28, not_a31b27, w_1_58_4, w_1_59_2);
	full_adder (not_a28b31, a29b30, a30b29, w_1_59_3, w_1_60_1);
	full_adder (not_a29b31, a30b30, not_a31b29, w_1_60_2, w_1_61_1);
	half_adder (not_a30b31, not_a31b30, w_1_61_2, w_1_62_1);
	half_adder (w_1_2_1, w_1_2_2, w_2_2_1, w_2_3_1);
	full_adder (w_1_3_1, w_1_3_2, a3b0, w_2_3_2, w_2_4_1);
	full_adder (w_1_4_1, w_1_4_2, w_1_4_3, w_2_4_2, w_2_5_1);
	full_adder (w_1_5_1, w_1_5_2, w_1_5_3, w_2_5_2, w_2_6_1);
	full_adder (w_1_6_1, w_1_6_2, w_1_6_3, w_2_6_2, w_2_7_1);
	half_adder (w_1_6_4, a6b0, w_2_6_3, w_2_7_2);
	full_adder (w_1_7_1, w_1_7_2, w_1_7_3, w_2_7_3, w_2_8_1);
	half_adder (w_1_7_4, w_1_7_5, w_2_7_4, w_2_8_2);
	full_adder (w_1_8_1, w_1_8_2, w_1_8_3, w_2_8_3, w_2_9_1);
	full_adder (w_1_8_4, w_1_8_5, w_1_8_6, w_2_8_4, w_2_9_2);
	full_adder (w_1_9_1, w_1_9_2, w_1_9_3, w_2_9_3, w_2_10_1);
	full_adder (w_1_9_4, w_1_9_5, w_1_9_6, w_2_9_4, w_2_10_2);
	full_adder (w_1_10_1, w_1_10_2, w_1_10_3, w_2_10_3, w_2_11_1);
	full_adder (w_1_10_4, w_1_10_5, w_1_10_6, w_2_10_4, w_2_11_2);
	full_adder (w_1_11_1, w_1_11_2, w_1_11_3, w_2_11_3, w_2_12_1);
	full_adder (w_1_11_4, w_1_11_5, w_1_11_6, w_2_11_4, w_2_12_2);
	half_adder (w_1_11_7, w_1_11_8, w_2_11_5, w_2_12_3);
	full_adder (w_1_12_1, w_1_12_2, w_1_12_3, w_2_12_4, w_2_13_1);
	full_adder (w_1_12_4, w_1_12_5, w_1_12_6, w_2_12_5, w_2_13_2);
	full_adder (w_1_12_7, w_1_12_8, a12b0, w_2_12_6, w_2_13_3);
	full_adder (w_1_13_1, w_1_13_2, w_1_13_3, w_2_13_4, w_2_14_1);
	full_adder (w_1_13_4, w_1_13_5, w_1_13_6, w_2_13_5, w_2_14_2);
	full_adder (w_1_13_7, w_1_13_8, w_1_13_9, w_2_13_6, w_2_14_3);
	full_adder (w_1_14_1, w_1_14_2, w_1_14_3, w_2_14_4, w_2_15_1);
	full_adder (w_1_14_4, w_1_14_5, w_1_14_6, w_2_14_5, w_2_15_2);
	full_adder (w_1_14_7, w_1_14_8, w_1_14_9, w_2_14_6, w_2_15_3);
	full_adder (w_1_15_1, w_1_15_2, w_1_15_3, w_2_15_4, w_2_16_1);
	full_adder (w_1_15_4, w_1_15_5, w_1_15_6, w_2_15_5, w_2_16_2);
	full_adder (w_1_15_7, w_1_15_8, w_1_15_9, w_2_15_6, w_2_16_3);
	half_adder (w_1_15_10, a15b0, w_2_15_7, w_2_16_4);
	full_adder (w_1_16_1, w_1_16_2, w_1_16_3, w_2_16_5, w_2_17_1);
	full_adder (w_1_16_4, w_1_16_5, w_1_16_6, w_2_16_6, w_2_17_2);
	full_adder (w_1_16_7, w_1_16_8, w_1_16_9, w_2_16_7, w_2_17_3);
	half_adder (w_1_16_10, w_1_16_11, w_2_16_8, w_2_17_4);
	full_adder (w_1_17_1, w_1_17_2, w_1_17_3, w_2_17_5, w_2_18_1);
	full_adder (w_1_17_4, w_1_17_5, w_1_17_6, w_2_17_6, w_2_18_2);
	full_adder (w_1_17_7, w_1_17_8, w_1_17_9, w_2_17_7, w_2_18_3);
	full_adder (w_1_17_10, w_1_17_11, w_1_17_12, w_2_17_8, w_2_18_4);
	full_adder (w_1_18_1, w_1_18_2, w_1_18_3, w_2_18_5, w_2_19_1);
	full_adder (w_1_18_4, w_1_18_5, w_1_18_6, w_2_18_6, w_2_19_2);
	full_adder (w_1_18_7, w_1_18_8, w_1_18_9, w_2_18_7, w_2_19_3);
	full_adder (w_1_18_10, w_1_18_11, w_1_18_12, w_2_18_8, w_2_19_4);
	full_adder (w_1_19_1, w_1_19_2, w_1_19_3, w_2_19_5, w_2_20_1);
	full_adder (w_1_19_4, w_1_19_5, w_1_19_6, w_2_19_6, w_2_20_2);
	full_adder (w_1_19_7, w_1_19_8, w_1_19_9, w_2_19_7, w_2_20_3);
	full_adder (w_1_19_10, w_1_19_11, w_1_19_12, w_2_19_8, w_2_20_4);
	full_adder (w_1_20_1, w_1_20_2, w_1_20_3, w_2_20_5, w_2_21_1);
	full_adder (w_1_20_4, w_1_20_5, w_1_20_6, w_2_20_6, w_2_21_2);
	full_adder (w_1_20_7, w_1_20_8, w_1_20_9, w_2_20_7, w_2_21_3);
	full_adder (w_1_20_10, w_1_20_11, w_1_20_12, w_2_20_8, w_2_21_4);
	half_adder (w_1_20_13, w_1_20_14, w_2_20_9, w_2_21_5);
	full_adder (w_1_21_1, w_1_21_2, w_1_21_3, w_2_21_6, w_2_22_1);
	full_adder (w_1_21_4, w_1_21_5, w_1_21_6, w_2_21_7, w_2_22_2);
	full_adder (w_1_21_7, w_1_21_8, w_1_21_9, w_2_21_8, w_2_22_3);
	full_adder (w_1_21_10, w_1_21_11, w_1_21_12, w_2_21_9, w_2_22_4);
	full_adder (w_1_21_13, w_1_21_14, a21b0, w_2_21_10, w_2_22_5);
	full_adder (w_1_22_1, w_1_22_2, w_1_22_3, w_2_22_6, w_2_23_1);
	full_adder (w_1_22_4, w_1_22_5, w_1_22_6, w_2_22_7, w_2_23_2);
	full_adder (w_1_22_7, w_1_22_8, w_1_22_9, w_2_22_8, w_2_23_3);
	full_adder (w_1_22_10, w_1_22_11, w_1_22_12, w_2_22_9, w_2_23_4);
	full_adder (w_1_22_13, w_1_22_14, w_1_22_15, w_2_22_10, w_2_23_5);
	full_adder (w_1_23_1, w_1_23_2, w_1_23_3, w_2_23_6, w_2_24_1);
	full_adder (w_1_23_4, w_1_23_5, w_1_23_6, w_2_23_7, w_2_24_2);
	full_adder (w_1_23_7, w_1_23_8, w_1_23_9, w_2_23_8, w_2_24_3);
	full_adder (w_1_23_10, w_1_23_11, w_1_23_12, w_2_23_9, w_2_24_4);
	full_adder (w_1_23_13, w_1_23_14, w_1_23_15, w_2_23_10, w_2_24_5);
	full_adder (w_1_24_1, w_1_24_2, w_1_24_3, w_2_24_6, w_2_25_1);
	full_adder (w_1_24_4, w_1_24_5, w_1_24_6, w_2_24_7, w_2_25_2);
	full_adder (w_1_24_7, w_1_24_8, w_1_24_9, w_2_24_8, w_2_25_3);
	full_adder (w_1_24_10, w_1_24_11, w_1_24_12, w_2_24_9, w_2_25_4);
	full_adder (w_1_24_13, w_1_24_14, w_1_24_15, w_2_24_10, w_2_25_5);
	half_adder (w_1_24_16, a24b0, w_2_24_11, w_2_25_6);
	full_adder (w_1_25_1, w_1_25_2, w_1_25_3, w_2_25_7, w_2_26_1);
	full_adder (w_1_25_4, w_1_25_5, w_1_25_6, w_2_25_8, w_2_26_2);
	full_adder (w_1_25_7, w_1_25_8, w_1_25_9, w_2_25_9, w_2_26_3);
	full_adder (w_1_25_10, w_1_25_11, w_1_25_12, w_2_25_10, w_2_26_4);
	full_adder (w_1_25_13, w_1_25_14, w_1_25_15, w_2_25_11, w_2_26_5);
	half_adder (w_1_25_16, w_1_25_17, w_2_25_12, w_2_26_6);
	full_adder (w_1_26_1, w_1_26_2, w_1_26_3, w_2_26_7, w_2_27_1);
	full_adder (w_1_26_4, w_1_26_5, w_1_26_6, w_2_26_8, w_2_27_2);
	full_adder (w_1_26_7, w_1_26_8, w_1_26_9, w_2_26_9, w_2_27_3);
	full_adder (w_1_26_10, w_1_26_11, w_1_26_12, w_2_26_10, w_2_27_4);
	full_adder (w_1_26_13, w_1_26_14, w_1_26_15, w_2_26_11, w_2_27_5);
	full_adder (w_1_26_16, w_1_26_17, w_1_26_18, w_2_26_12, w_2_27_6);
	full_adder (w_1_27_1, w_1_27_2, w_1_27_3, w_2_27_7, w_2_28_1);
	full_adder (w_1_27_4, w_1_27_5, w_1_27_6, w_2_27_8, w_2_28_2);
	full_adder (w_1_27_7, w_1_27_8, w_1_27_9, w_2_27_9, w_2_28_3);
	full_adder (w_1_27_10, w_1_27_11, w_1_27_12, w_2_27_10, w_2_28_4);
	full_adder (w_1_27_13, w_1_27_14, w_1_27_15, w_2_27_11, w_2_28_5);
	full_adder (w_1_27_16, w_1_27_17, w_1_27_18, w_2_27_12, w_2_28_6);
	full_adder (w_1_28_1, w_1_28_2, w_1_28_3, w_2_28_7, w_2_29_1);
	full_adder (w_1_28_4, w_1_28_5, w_1_28_6, w_2_28_8, w_2_29_2);
	full_adder (w_1_28_7, w_1_28_8, w_1_28_9, w_2_28_9, w_2_29_3);
	full_adder (w_1_28_10, w_1_28_11, w_1_28_12, w_2_28_10, w_2_29_4);
	full_adder (w_1_28_13, w_1_28_14, w_1_28_15, w_2_28_11, w_2_29_5);
	full_adder (w_1_28_16, w_1_28_17, w_1_28_18, w_2_28_12, w_2_29_6);
	full_adder (w_1_29_1, w_1_29_2, w_1_29_3, w_2_29_7, w_2_30_1);
	full_adder (w_1_29_4, w_1_29_5, w_1_29_6, w_2_29_8, w_2_30_2);
	full_adder (w_1_29_7, w_1_29_8, w_1_29_9, w_2_29_9, w_2_30_3);
	full_adder (w_1_29_10, w_1_29_11, w_1_29_12, w_2_29_10, w_2_30_4);
	full_adder (w_1_29_13, w_1_29_14, w_1_29_15, w_2_29_11, w_2_30_5);
	full_adder (w_1_29_16, w_1_29_17, w_1_29_18, w_2_29_12, w_2_30_6);
	half_adder (w_1_29_19, w_1_29_20, w_2_29_13, w_2_30_7);
	full_adder (w_1_30_1, w_1_30_2, w_1_30_3, w_2_30_8, w_2_31_1);
	full_adder (w_1_30_4, w_1_30_5, w_1_30_6, w_2_30_9, w_2_31_2);
	full_adder (w_1_30_7, w_1_30_8, w_1_30_9, w_2_30_10, w_2_31_3);
	full_adder (w_1_30_10, w_1_30_11, w_1_30_12, w_2_30_11, w_2_31_4);
	full_adder (w_1_30_13, w_1_30_14, w_1_30_15, w_2_30_12, w_2_31_5);
	full_adder (w_1_30_16, w_1_30_17, w_1_30_18, w_2_30_13, w_2_31_6);
	full_adder (w_1_30_19, w_1_30_20, a30b0, w_2_30_14, w_2_31_7);
	full_adder (w_1_31_1, w_1_31_2, w_1_31_3, w_2_31_8, w_2_32_1);
	full_adder (w_1_31_4, w_1_31_5, w_1_31_6, w_2_31_9, w_2_32_2);
	full_adder (w_1_31_7, w_1_31_8, w_1_31_9, w_2_31_10, w_2_32_3);
	full_adder (w_1_31_10, w_1_31_11, w_1_31_12, w_2_31_11, w_2_32_4);
	full_adder (w_1_31_13, w_1_31_14, w_1_31_15, w_2_31_12, w_2_32_5);
	full_adder (w_1_31_16, w_1_31_17, w_1_31_18, w_2_31_13, w_2_32_6);
	full_adder (w_1_31_19, w_1_31_20, w_1_31_21, w_2_31_14, w_2_32_7);
	full_adder (w_1_32_1, w_1_32_2, w_1_32_3, w_2_32_8, w_2_33_1);
	full_adder (w_1_32_4, w_1_32_5, w_1_32_6, w_2_32_9, w_2_33_2);
	full_adder (w_1_32_7, w_1_32_8, w_1_32_9, w_2_32_10, w_2_33_3);
	full_adder (w_1_32_10, w_1_32_11, w_1_32_12, w_2_32_11, w_2_33_4);
	full_adder (w_1_32_13, w_1_32_14, w_1_32_15, w_2_32_12, w_2_33_5);
	full_adder (w_1_32_16, w_1_32_17, w_1_32_18, w_2_32_13, w_2_33_6);
	full_adder (w_1_32_19, w_1_32_20, w_1_32_21, w_2_32_14, w_2_33_7);
	full_adder (w_1_33_1, w_1_33_2, w_1_33_3, w_2_33_8, w_2_34_1);
	full_adder (w_1_33_4, w_1_33_5, w_1_33_6, w_2_33_9, w_2_34_2);
	full_adder (w_1_33_7, w_1_33_8, w_1_33_9, w_2_33_10, w_2_34_3);
	full_adder (w_1_33_10, w_1_33_11, w_1_33_12, w_2_33_11, w_2_34_4);
	full_adder (w_1_33_13, w_1_33_14, w_1_33_15, w_2_33_12, w_2_34_5);
	full_adder (w_1_33_16, w_1_33_17, w_1_33_18, w_2_33_13, w_2_34_6);
	full_adder (w_1_33_19, w_1_33_20, w_1_33_21, w_2_33_14, w_2_34_7);
	full_adder (w_1_34_1, w_1_34_2, w_1_34_3, w_2_34_8, w_2_35_1);
	full_adder (w_1_34_4, w_1_34_5, w_1_34_6, w_2_34_9, w_2_35_2);
	full_adder (w_1_34_7, w_1_34_8, w_1_34_9, w_2_34_10, w_2_35_3);
	full_adder (w_1_34_10, w_1_34_11, w_1_34_12, w_2_34_11, w_2_35_4);
	full_adder (w_1_34_13, w_1_34_14, w_1_34_15, w_2_34_12, w_2_35_5);
	full_adder (w_1_34_16, w_1_34_17, w_1_34_18, w_2_34_13, w_2_35_6);
	half_adder (w_1_34_19, w_1_34_20, w_2_34_14, w_2_35_7);
	full_adder (w_1_35_1, w_1_35_2, w_1_35_3, w_2_35_8, w_2_36_1);
	full_adder (w_1_35_4, w_1_35_5, w_1_35_6, w_2_35_9, w_2_36_2);
	full_adder (w_1_35_7, w_1_35_8, w_1_35_9, w_2_35_10, w_2_36_3);
	full_adder (w_1_35_10, w_1_35_11, w_1_35_12, w_2_35_11, w_2_36_4);
	full_adder (w_1_35_13, w_1_35_14, w_1_35_15, w_2_35_12, w_2_36_5);
	full_adder (w_1_35_16, w_1_35_17, w_1_35_18, w_2_35_13, w_2_36_6);
	half_adder (w_1_35_19, not_a31b4, w_2_35_14, w_2_36_7);
	full_adder (w_1_36_1, w_1_36_2, w_1_36_3, w_2_36_8, w_2_37_1);
	full_adder (w_1_36_4, w_1_36_5, w_1_36_6, w_2_36_9, w_2_37_2);
	full_adder (w_1_36_7, w_1_36_8, w_1_36_9, w_2_36_10, w_2_37_3);
	full_adder (w_1_36_10, w_1_36_11, w_1_36_12, w_2_36_11, w_2_37_4);
	full_adder (w_1_36_13, w_1_36_14, w_1_36_15, w_2_36_12, w_2_37_5);
	full_adder (w_1_36_16, w_1_36_17, w_1_36_18, w_2_36_13, w_2_37_6);
	full_adder (w_1_37_1, w_1_37_2, w_1_37_3, w_2_37_7, w_2_38_1);
	full_adder (w_1_37_4, w_1_37_5, w_1_37_6, w_2_37_8, w_2_38_2);
	full_adder (w_1_37_7, w_1_37_8, w_1_37_9, w_2_37_9, w_2_38_3);
	full_adder (w_1_37_10, w_1_37_11, w_1_37_12, w_2_37_10, w_2_38_4);
	full_adder (w_1_37_13, w_1_37_14, w_1_37_15, w_2_37_11, w_2_38_5);
	full_adder (w_1_37_16, w_1_37_17, w_1_37_18, w_2_37_12, w_2_38_6);
	full_adder (w_1_38_1, w_1_38_2, w_1_38_3, w_2_38_7, w_2_39_1);
	full_adder (w_1_38_4, w_1_38_5, w_1_38_6, w_2_38_8, w_2_39_2);
	full_adder (w_1_38_7, w_1_38_8, w_1_38_9, w_2_38_9, w_2_39_3);
	full_adder (w_1_38_10, w_1_38_11, w_1_38_12, w_2_38_10, w_2_39_4);
	full_adder (w_1_38_13, w_1_38_14, w_1_38_15, w_2_38_11, w_2_39_5);
	full_adder (w_1_38_16, w_1_38_17, not_a31b7, w_2_38_12, w_2_39_6);
	full_adder (w_1_39_1, w_1_39_2, w_1_39_3, w_2_39_7, w_2_40_1);
	full_adder (w_1_39_4, w_1_39_5, w_1_39_6, w_2_39_8, w_2_40_2);
	full_adder (w_1_39_7, w_1_39_8, w_1_39_9, w_2_39_9, w_2_40_3);
	full_adder (w_1_39_10, w_1_39_11, w_1_39_12, w_2_39_10, w_2_40_4);
	full_adder (w_1_39_13, w_1_39_14, w_1_39_15, w_2_39_11, w_2_40_5);
	full_adder (w_1_40_1, w_1_40_2, w_1_40_3, w_2_40_6, w_2_41_1);
	full_adder (w_1_40_4, w_1_40_5, w_1_40_6, w_2_40_7, w_2_41_2);
	full_adder (w_1_40_7, w_1_40_8, w_1_40_9, w_2_40_8, w_2_41_3);
	full_adder (w_1_40_10, w_1_40_11, w_1_40_12, w_2_40_9, w_2_41_4);
	full_adder (w_1_40_13, w_1_40_14, w_1_40_15, w_2_40_10, w_2_41_5);
	full_adder (w_1_41_1, w_1_41_2, w_1_41_3, w_2_41_6, w_2_42_1);
	full_adder (w_1_41_4, w_1_41_5, w_1_41_6, w_2_41_7, w_2_42_2);
	full_adder (w_1_41_7, w_1_41_8, w_1_41_9, w_2_41_8, w_2_42_3);
	full_adder (w_1_41_10, w_1_41_11, w_1_41_12, w_2_41_9, w_2_42_4);
	full_adder (w_1_41_13, w_1_41_14, w_1_41_15, w_2_41_10, w_2_42_5);
	full_adder (w_1_42_1, w_1_42_2, w_1_42_3, w_2_42_6, w_2_43_1);
	full_adder (w_1_42_4, w_1_42_5, w_1_42_6, w_2_42_7, w_2_43_2);
	full_adder (w_1_42_7, w_1_42_8, w_1_42_9, w_2_42_8, w_2_43_3);
	full_adder (w_1_42_10, w_1_42_11, w_1_42_12, w_2_42_9, w_2_43_4);
	half_adder (w_1_42_13, w_1_42_14, w_2_42_10, w_2_43_5);
	full_adder (w_1_43_1, w_1_43_2, w_1_43_3, w_2_43_6, w_2_44_1);
	full_adder (w_1_43_4, w_1_43_5, w_1_43_6, w_2_43_7, w_2_44_2);
	full_adder (w_1_43_7, w_1_43_8, w_1_43_9, w_2_43_8, w_2_44_3);
	full_adder (w_1_43_10, w_1_43_11, w_1_43_12, w_2_43_9, w_2_44_4);
	half_adder (w_1_43_13, w_1_43_14, w_2_43_10, w_2_44_5);
	full_adder (w_1_44_1, w_1_44_2, w_1_44_3, w_2_44_6, w_2_45_1);
	full_adder (w_1_44_4, w_1_44_5, w_1_44_6, w_2_44_7, w_2_45_2);
	full_adder (w_1_44_7, w_1_44_8, w_1_44_9, w_2_44_8, w_2_45_3);
	full_adder (w_1_44_10, w_1_44_11, w_1_44_12, w_2_44_9, w_2_45_4);
	half_adder (w_1_44_13, not_a31b13, w_2_44_10, w_2_45_5);
	full_adder (w_1_45_1, w_1_45_2, w_1_45_3, w_2_45_6, w_2_46_1);
	full_adder (w_1_45_4, w_1_45_5, w_1_45_6, w_2_45_7, w_2_46_2);
	full_adder (w_1_45_7, w_1_45_8, w_1_45_9, w_2_45_8, w_2_46_3);
	full_adder (w_1_45_10, w_1_45_11, w_1_45_12, w_2_45_9, w_2_46_4);
	full_adder (w_1_46_1, w_1_46_2, w_1_46_3, w_2_46_5, w_2_47_1);
	full_adder (w_1_46_4, w_1_46_5, w_1_46_6, w_2_46_6, w_2_47_2);
	full_adder (w_1_46_7, w_1_46_8, w_1_46_9, w_2_46_7, w_2_47_3);
	full_adder (w_1_46_10, w_1_46_11, w_1_46_12, w_2_46_8, w_2_47_4);
	full_adder (w_1_47_1, w_1_47_2, w_1_47_3, w_2_47_5, w_2_48_1);
	full_adder (w_1_47_4, w_1_47_5, w_1_47_6, w_2_47_6, w_2_48_2);
	full_adder (w_1_47_7, w_1_47_8, w_1_47_9, w_2_47_7, w_2_48_3);
	full_adder (w_1_47_10, w_1_47_11, not_a31b16, w_2_47_8, w_2_48_4);
	full_adder (w_1_48_1, w_1_48_2, w_1_48_3, w_2_48_5, w_2_49_1);
	full_adder (w_1_48_4, w_1_48_5, w_1_48_6, w_2_48_6, w_2_49_2);
	full_adder (w_1_48_7, w_1_48_8, w_1_48_9, w_2_48_7, w_2_49_3);
	full_adder (w_1_49_1, w_1_49_2, w_1_49_3, w_2_49_4, w_2_50_1);
	full_adder (w_1_49_4, w_1_49_5, w_1_49_6, w_2_49_5, w_2_50_2);
	full_adder (w_1_49_7, w_1_49_8, w_1_49_9, w_2_49_6, w_2_50_3);
	full_adder (w_1_50_1, w_1_50_2, w_1_50_3, w_2_50_4, w_2_51_1);
	full_adder (w_1_50_4, w_1_50_5, w_1_50_6, w_2_50_5, w_2_51_2);
	full_adder (w_1_50_7, w_1_50_8, w_1_50_9, w_2_50_6, w_2_51_3);
	full_adder (w_1_51_1, w_1_51_2, w_1_51_3, w_2_51_4, w_2_52_1);
	full_adder (w_1_51_4, w_1_51_5, w_1_51_6, w_2_51_5, w_2_52_2);
	half_adder (w_1_51_7, w_1_51_8, w_2_51_6, w_2_52_3);
	full_adder (w_1_52_1, w_1_52_2, w_1_52_3, w_2_52_4, w_2_53_1);
	full_adder (w_1_52_4, w_1_52_5, w_1_52_6, w_2_52_5, w_2_53_2);
	half_adder (w_1_52_7, w_1_52_8, w_2_52_6, w_2_53_3);
	full_adder (w_1_53_1, w_1_53_2, w_1_53_3, w_2_53_4, w_2_54_1);
	full_adder (w_1_53_4, w_1_53_5, w_1_53_6, w_2_53_5, w_2_54_2);
	half_adder (w_1_53_7, not_a31b22, w_2_53_6, w_2_54_3);
	full_adder (w_1_54_1, w_1_54_2, w_1_54_3, w_2_54_4, w_2_55_1);
	full_adder (w_1_54_4, w_1_54_5, w_1_54_6, w_2_54_5, w_2_55_2);
	full_adder (w_1_55_1, w_1_55_2, w_1_55_3, w_2_55_3, w_2_56_1);
	full_adder (w_1_55_4, w_1_55_5, w_1_55_6, w_2_55_4, w_2_56_2);
	full_adder (w_1_56_1, w_1_56_2, w_1_56_3, w_2_56_3, w_2_57_1);
	full_adder (w_1_56_4, w_1_56_5, not_a31b25, w_2_56_4, w_2_57_2);
	full_adder (w_1_57_1, w_1_57_2, w_1_57_3, w_2_57_3, w_2_58_1);
	full_adder (w_1_58_1, w_1_58_2, w_1_58_3, w_2_58_2, w_2_59_1);
	full_adder (w_1_59_1, w_1_59_2, w_1_59_3, w_2_59_2, w_2_60_1);
	half_adder (w_1_60_1, w_1_60_2, w_2_60_2, w_2_61_1);
	half_adder (w_1_61_1, w_1_61_2, w_2_61_2, w_2_62_1);
	half_adder (w_1_62_1, a31b31, w_2_62_2, w_2_63_1);
	half_adder (w_2_3_1, w_2_3_2, w_3_3_1, w_3_4_1);
	half_adder (w_2_4_1, w_2_4_2, w_3_4_2, w_3_5_1);
	full_adder (w_2_5_1, w_2_5_2, w_1_5_4, w_3_5_2, w_3_6_1);
	full_adder (w_2_6_1, w_2_6_2, w_2_6_3, w_3_6_2, w_3_7_1);
	full_adder (w_2_7_1, w_2_7_2, w_2_7_3, w_3_7_2, w_3_8_1);
	full_adder (w_2_8_1, w_2_8_2, w_2_8_3, w_3_8_2, w_3_9_1);
	full_adder (w_2_9_1, w_2_9_2, w_2_9_3, w_3_9_2, w_3_10_1);
	half_adder (w_2_9_4, a9b0, w_3_9_3, w_3_10_2);
	full_adder (w_2_10_1, w_2_10_2, w_2_10_3, w_3_10_3, w_3_11_1);
	half_adder (w_2_10_4, w_1_10_7, w_3_10_4, w_3_11_2);
	full_adder (w_2_11_1, w_2_11_2, w_2_11_3, w_3_11_3, w_3_12_1);
	half_adder (w_2_11_4, w_2_11_5, w_3_11_4, w_3_12_2);
	full_adder (w_2_12_1, w_2_12_2, w_2_12_3, w_3_12_3, w_3_13_1);
	full_adder (w_2_12_4, w_2_12_5, w_2_12_6, w_3_12_4, w_3_13_2);
	full_adder (w_2_13_1, w_2_13_2, w_2_13_3, w_3_13_3, w_3_14_1);
	full_adder (w_2_13_4, w_2_13_5, w_2_13_6, w_3_13_4, w_3_14_2);
	full_adder (w_2_14_1, w_2_14_2, w_2_14_3, w_3_14_3, w_3_15_1);
	full_adder (w_2_14_4, w_2_14_5, w_2_14_6, w_3_14_4, w_3_15_2);
	full_adder (w_2_15_1, w_2_15_2, w_2_15_3, w_3_15_3, w_3_16_1);
	full_adder (w_2_15_4, w_2_15_5, w_2_15_6, w_3_15_4, w_3_16_2);
	full_adder (w_2_16_1, w_2_16_2, w_2_16_3, w_3_16_3, w_3_17_1);
	full_adder (w_2_16_4, w_2_16_5, w_2_16_6, w_3_16_4, w_3_17_2);
	half_adder (w_2_16_7, w_2_16_8, w_3_16_5, w_3_17_3);
	full_adder (w_2_17_1, w_2_17_2, w_2_17_3, w_3_17_4, w_3_18_1);
	full_adder (w_2_17_4, w_2_17_5, w_2_17_6, w_3_17_5, w_3_18_2);
	half_adder (w_2_17_7, w_2_17_8, w_3_17_6, w_3_18_3);
	full_adder (w_2_18_1, w_2_18_2, w_2_18_3, w_3_18_4, w_3_19_1);
	full_adder (w_2_18_4, w_2_18_5, w_2_18_6, w_3_18_5, w_3_19_2);
	full_adder (w_2_18_7, w_2_18_8, a18b0, w_3_18_6, w_3_19_3);
	full_adder (w_2_19_1, w_2_19_2, w_2_19_3, w_3_19_4, w_3_20_1);
	full_adder (w_2_19_4, w_2_19_5, w_2_19_6, w_3_19_5, w_3_20_2);
	full_adder (w_2_19_7, w_2_19_8, w_1_19_13, w_3_19_6, w_3_20_3);
	full_adder (w_2_20_1, w_2_20_2, w_2_20_3, w_3_20_4, w_3_21_1);
	full_adder (w_2_20_4, w_2_20_5, w_2_20_6, w_3_20_5, w_3_21_2);
	full_adder (w_2_20_7, w_2_20_8, w_2_20_9, w_3_20_6, w_3_21_3);
	full_adder (w_2_21_1, w_2_21_2, w_2_21_3, w_3_21_4, w_3_22_1);
	full_adder (w_2_21_4, w_2_21_5, w_2_21_6, w_3_21_5, w_3_22_2);
	full_adder (w_2_21_7, w_2_21_8, w_2_21_9, w_3_21_6, w_3_22_3);
	full_adder (w_2_22_1, w_2_22_2, w_2_22_3, w_3_22_4, w_3_23_1);
	full_adder (w_2_22_4, w_2_22_5, w_2_22_6, w_3_22_5, w_3_23_2);
	full_adder (w_2_22_7, w_2_22_8, w_2_22_9, w_3_22_6, w_3_23_3);
	full_adder (w_2_23_1, w_2_23_2, w_2_23_3, w_3_23_4, w_3_24_1);
	full_adder (w_2_23_4, w_2_23_5, w_2_23_6, w_3_23_5, w_3_24_2);
	full_adder (w_2_23_7, w_2_23_8, w_2_23_9, w_3_23_6, w_3_24_3);
	half_adder (w_2_23_10, w_1_23_16, w_3_23_7, w_3_24_4);
	full_adder (w_2_24_1, w_2_24_2, w_2_24_3, w_3_24_5, w_3_25_1);
	full_adder (w_2_24_4, w_2_24_5, w_2_24_6, w_3_24_6, w_3_25_2);
	full_adder (w_2_24_7, w_2_24_8, w_2_24_9, w_3_24_7, w_3_25_3);
	half_adder (w_2_24_10, w_2_24_11, w_3_24_8, w_3_25_4);
	full_adder (w_2_25_1, w_2_25_2, w_2_25_3, w_3_25_5, w_3_26_1);
	full_adder (w_2_25_4, w_2_25_5, w_2_25_6, w_3_25_6, w_3_26_2);
	full_adder (w_2_25_7, w_2_25_8, w_2_25_9, w_3_25_7, w_3_26_3);
	full_adder (w_2_25_10, w_2_25_11, w_2_25_12, w_3_25_8, w_3_26_4);
	full_adder (w_2_26_1, w_2_26_2, w_2_26_3, w_3_26_5, w_3_27_1);
	full_adder (w_2_26_4, w_2_26_5, w_2_26_6, w_3_26_6, w_3_27_2);
	full_adder (w_2_26_7, w_2_26_8, w_2_26_9, w_3_26_7, w_3_27_3);
	full_adder (w_2_26_10, w_2_26_11, w_2_26_12, w_3_26_8, w_3_27_4);
	full_adder (w_2_27_1, w_2_27_2, w_2_27_3, w_3_27_5, w_3_28_1);
	full_adder (w_2_27_4, w_2_27_5, w_2_27_6, w_3_27_6, w_3_28_2);
	full_adder (w_2_27_7, w_2_27_8, w_2_27_9, w_3_27_7, w_3_28_3);
	full_adder (w_2_27_10, w_2_27_11, w_2_27_12, w_3_27_8, w_3_28_4);
	full_adder (w_2_28_1, w_2_28_2, w_2_28_3, w_3_28_5, w_3_29_1);
	full_adder (w_2_28_4, w_2_28_5, w_2_28_6, w_3_28_6, w_3_29_2);
	full_adder (w_2_28_7, w_2_28_8, w_2_28_9, w_3_28_7, w_3_29_3);
	full_adder (w_2_28_10, w_2_28_11, w_2_28_12, w_3_28_8, w_3_29_4);
	full_adder (w_2_29_1, w_2_29_2, w_2_29_3, w_3_29_5, w_3_30_1);
	full_adder (w_2_29_4, w_2_29_5, w_2_29_6, w_3_29_6, w_3_30_2);
	full_adder (w_2_29_7, w_2_29_8, w_2_29_9, w_3_29_7, w_3_30_3);
	full_adder (w_2_29_10, w_2_29_11, w_2_29_12, w_3_29_8, w_3_30_4);
	full_adder (w_2_30_1, w_2_30_2, w_2_30_3, w_3_30_5, w_3_31_1);
	full_adder (w_2_30_4, w_2_30_5, w_2_30_6, w_3_30_6, w_3_31_2);
	full_adder (w_2_30_7, w_2_30_8, w_2_30_9, w_3_30_7, w_3_31_3);
	full_adder (w_2_30_10, w_2_30_11, w_2_30_12, w_3_30_8, w_3_31_4);
	half_adder (w_2_30_13, w_2_30_14, w_3_30_9, w_3_31_5);
	full_adder (w_2_31_1, w_2_31_2, w_2_31_3, w_3_31_6, w_3_32_1);
	full_adder (w_2_31_4, w_2_31_5, w_2_31_6, w_3_31_7, w_3_32_2);
	full_adder (w_2_31_7, w_2_31_8, w_2_31_9, w_3_31_8, w_3_32_3);
	full_adder (w_2_31_10, w_2_31_11, w_2_31_12, w_3_31_9, w_3_32_4);
	half_adder (w_2_31_13, w_2_31_14, w_3_31_10, w_3_32_5);
	full_adder (w_2_32_1, w_2_32_2, w_2_32_3, w_3_32_6, w_3_33_1);
	full_adder (w_2_32_4, w_2_32_5, w_2_32_6, w_3_32_7, w_3_33_2);
	full_adder (w_2_32_7, w_2_32_8, w_2_32_9, w_3_32_8, w_3_33_3);
	full_adder (w_2_32_10, w_2_32_11, w_2_32_12, w_3_32_9, w_3_33_4);
	full_adder (w_2_32_13, w_2_32_14, w_1_32_22, w_3_32_10, w_3_33_5);
	full_adder (w_2_33_1, w_2_33_2, w_2_33_3, w_3_33_6, w_3_34_1);
	full_adder (w_2_33_4, w_2_33_5, w_2_33_6, w_3_33_7, w_3_34_2);
	full_adder (w_2_33_7, w_2_33_8, w_2_33_9, w_3_33_8, w_3_34_3);
	full_adder (w_2_33_10, w_2_33_11, w_2_33_12, w_3_33_9, w_3_34_4);
	half_adder (w_2_33_13, w_2_33_14, w_3_33_10, w_3_34_5);
	full_adder (w_2_34_1, w_2_34_2, w_2_34_3, w_3_34_6, w_3_35_1);
	full_adder (w_2_34_4, w_2_34_5, w_2_34_6, w_3_34_7, w_3_35_2);
	full_adder (w_2_34_7, w_2_34_8, w_2_34_9, w_3_34_8, w_3_35_3);
	full_adder (w_2_34_10, w_2_34_11, w_2_34_12, w_3_34_9, w_3_35_4);
	half_adder (w_2_34_13, w_2_34_14, w_3_34_10, w_3_35_5);
	full_adder (w_2_35_1, w_2_35_2, w_2_35_3, w_3_35_6, w_3_36_1);
	full_adder (w_2_35_4, w_2_35_5, w_2_35_6, w_3_35_7, w_3_36_2);
	full_adder (w_2_35_7, w_2_35_8, w_2_35_9, w_3_35_8, w_3_36_3);
	full_adder (w_2_35_10, w_2_35_11, w_2_35_12, w_3_35_9, w_3_36_4);
	half_adder (w_2_35_13, w_2_35_14, w_3_35_10, w_3_36_5);
	full_adder (w_2_36_1, w_2_36_2, w_2_36_3, w_3_36_6, w_3_37_1);
	full_adder (w_2_36_4, w_2_36_5, w_2_36_6, w_3_36_7, w_3_37_2);
	full_adder (w_2_36_7, w_2_36_8, w_2_36_9, w_3_36_8, w_3_37_3);
	full_adder (w_2_36_10, w_2_36_11, w_2_36_12, w_3_36_9, w_3_37_4);
	full_adder (w_2_37_1, w_2_37_2, w_2_37_3, w_3_37_5, w_3_38_1);
	full_adder (w_2_37_4, w_2_37_5, w_2_37_6, w_3_37_6, w_3_38_2);
	full_adder (w_2_37_7, w_2_37_8, w_2_37_9, w_3_37_7, w_3_38_3);
	full_adder (w_2_37_10, w_2_37_11, w_2_37_12, w_3_37_8, w_3_38_4);
	full_adder (w_2_38_1, w_2_38_2, w_2_38_3, w_3_38_5, w_3_39_1);
	full_adder (w_2_38_4, w_2_38_5, w_2_38_6, w_3_38_6, w_3_39_2);
	full_adder (w_2_38_7, w_2_38_8, w_2_38_9, w_3_38_7, w_3_39_3);
	full_adder (w_2_38_10, w_2_38_11, w_2_38_12, w_3_38_8, w_3_39_4);
	full_adder (w_2_39_1, w_2_39_2, w_2_39_3, w_3_39_5, w_3_40_1);
	full_adder (w_2_39_4, w_2_39_5, w_2_39_6, w_3_39_6, w_3_40_2);
	full_adder (w_2_39_7, w_2_39_8, w_2_39_9, w_3_39_7, w_3_40_3);
	full_adder (w_2_39_10, w_2_39_11, w_1_39_16, w_3_39_8, w_3_40_4);
	full_adder (w_2_40_1, w_2_40_2, w_2_40_3, w_3_40_5, w_3_41_1);
	full_adder (w_2_40_4, w_2_40_5, w_2_40_6, w_3_40_6, w_3_41_2);
	full_adder (w_2_40_7, w_2_40_8, w_2_40_9, w_3_40_7, w_3_41_3);
	half_adder (w_2_40_10, w_1_40_16, w_3_40_8, w_3_41_4);
	full_adder (w_2_41_1, w_2_41_2, w_2_41_3, w_3_41_5, w_3_42_1);
	full_adder (w_2_41_4, w_2_41_5, w_2_41_6, w_3_41_6, w_3_42_2);
	full_adder (w_2_41_7, w_2_41_8, w_2_41_9, w_3_41_7, w_3_42_3);
	half_adder (w_2_41_10, not_a31b10, w_3_41_8, w_3_42_4);
	full_adder (w_2_42_1, w_2_42_2, w_2_42_3, w_3_42_5, w_3_43_1);
	full_adder (w_2_42_4, w_2_42_5, w_2_42_6, w_3_42_6, w_3_43_2);
	full_adder (w_2_42_7, w_2_42_8, w_2_42_9, w_3_42_7, w_3_43_3);
	full_adder (w_2_43_1, w_2_43_2, w_2_43_3, w_3_43_4, w_3_44_1);
	full_adder (w_2_43_4, w_2_43_5, w_2_43_6, w_3_43_5, w_3_44_2);
	full_adder (w_2_43_7, w_2_43_8, w_2_43_9, w_3_43_6, w_3_44_3);
	full_adder (w_2_44_1, w_2_44_2, w_2_44_3, w_3_44_4, w_3_45_1);
	full_adder (w_2_44_4, w_2_44_5, w_2_44_6, w_3_44_5, w_3_45_2);
	full_adder (w_2_44_7, w_2_44_8, w_2_44_9, w_3_44_6, w_3_45_3);
	full_adder (w_2_45_1, w_2_45_2, w_2_45_3, w_3_45_4, w_3_46_1);
	full_adder (w_2_45_4, w_2_45_5, w_2_45_6, w_3_45_5, w_3_46_2);
	full_adder (w_2_45_7, w_2_45_8, w_2_45_9, w_3_45_6, w_3_46_3);
	full_adder (w_2_46_1, w_2_46_2, w_2_46_3, w_3_46_4, w_3_47_1);
	full_adder (w_2_46_4, w_2_46_5, w_2_46_6, w_3_46_5, w_3_47_2);
	half_adder (w_2_46_7, w_2_46_8, w_3_46_6, w_3_47_3);
	full_adder (w_2_47_1, w_2_47_2, w_2_47_3, w_3_47_4, w_3_48_1);
	full_adder (w_2_47_4, w_2_47_5, w_2_47_6, w_3_47_5, w_3_48_2);
	half_adder (w_2_47_7, w_2_47_8, w_3_47_6, w_3_48_3);
	full_adder (w_2_48_1, w_2_48_2, w_2_48_3, w_3_48_4, w_3_49_1);
	full_adder (w_2_48_4, w_2_48_5, w_2_48_6, w_3_48_5, w_3_49_2);
	half_adder (w_2_48_7, w_1_48_10, w_3_48_6, w_3_49_3);
	full_adder (w_2_49_1, w_2_49_2, w_2_49_3, w_3_49_4, w_3_50_1);
	full_adder (w_2_49_4, w_2_49_5, w_2_49_6, w_3_49_5, w_3_50_2);
	full_adder (w_2_50_1, w_2_50_2, w_2_50_3, w_3_50_3, w_3_51_1);
	full_adder (w_2_50_4, w_2_50_5, w_2_50_6, w_3_50_4, w_3_51_2);
	full_adder (w_2_51_1, w_2_51_2, w_2_51_3, w_3_51_3, w_3_52_1);
	full_adder (w_2_51_4, w_2_51_5, w_2_51_6, w_3_51_4, w_3_52_2);
	full_adder (w_2_52_1, w_2_52_2, w_2_52_3, w_3_52_3, w_3_53_1);
	full_adder (w_2_52_4, w_2_52_5, w_2_52_6, w_3_52_4, w_3_53_2);
	full_adder (w_2_53_1, w_2_53_2, w_2_53_3, w_3_53_3, w_3_54_1);
	full_adder (w_2_53_4, w_2_53_5, w_2_53_6, w_3_53_4, w_3_54_2);
	full_adder (w_2_54_1, w_2_54_2, w_2_54_3, w_3_54_3, w_3_55_1);
	half_adder (w_2_54_4, w_2_54_5, w_3_54_4, w_3_55_2);
	full_adder (w_2_55_1, w_2_55_2, w_2_55_3, w_3_55_3, w_3_56_1);
	full_adder (w_2_56_1, w_2_56_2, w_2_56_3, w_3_56_2, w_3_57_1);
	full_adder (w_2_57_1, w_2_57_2, w_2_57_3, w_3_57_2, w_3_58_1);
	full_adder (w_2_58_1, w_2_58_2, w_1_58_4, w_3_58_2, w_3_59_1);
	full_adder (w_2_59_1, w_2_59_2, not_a31b28, w_3_59_2, w_3_60_1);
	half_adder (w_2_60_1, w_2_60_2, w_3_60_2, w_3_61_1);
	half_adder (w_2_61_1, w_2_61_2, w_3_61_2, w_3_62_1);
	half_adder (w_2_62_1, w_2_62_2, w_3_62_2, w_3_63_1);
	half_adder (w_2_63_1, 1, w_3_63_2, w_3_64_1);
	half_adder (w_3_4_1, w_3_4_2, w_4_4_1, w_4_5_1);
	half_adder (w_3_5_1, w_3_5_2, w_4_5_2, w_4_6_1);
	half_adder (w_3_6_1, w_3_6_2, w_4_6_2, w_4_7_1);
	full_adder (w_3_7_1, w_3_7_2, w_2_7_4, w_4_7_2, w_4_8_1);
	full_adder (w_3_8_1, w_3_8_2, w_2_8_4, w_4_8_2, w_4_9_1);
	full_adder (w_3_9_1, w_3_9_2, w_3_9_3, w_4_9_2, w_4_10_1);
	full_adder (w_3_10_1, w_3_10_2, w_3_10_3, w_4_10_2, w_4_11_1);
	full_adder (w_3_11_1, w_3_11_2, w_3_11_3, w_4_11_2, w_4_12_1);
	full_adder (w_3_12_1, w_3_12_2, w_3_12_3, w_4_12_2, w_4_13_1);
	full_adder (w_3_13_1, w_3_13_2, w_3_13_3, w_4_13_2, w_4_14_1);
	full_adder (w_3_14_1, w_3_14_2, w_3_14_3, w_4_14_2, w_4_15_1);
	half_adder (w_3_14_4, w_1_14_10, w_4_14_3, w_4_15_2);
	full_adder (w_3_15_1, w_3_15_2, w_3_15_3, w_4_15_3, w_4_16_1);
	half_adder (w_3_15_4, w_2_15_7, w_4_15_4, w_4_16_2);
	full_adder (w_3_16_1, w_3_16_2, w_3_16_3, w_4_16_3, w_4_17_1);
	half_adder (w_3_16_4, w_3_16_5, w_4_16_4, w_4_17_2);
	full_adder (w_3_17_1, w_3_17_2, w_3_17_3, w_4_17_3, w_4_18_1);
	full_adder (w_3_17_4, w_3_17_5, w_3_17_6, w_4_17_4, w_4_18_2);
	full_adder (w_3_18_1, w_3_18_2, w_3_18_3, w_4_18_3, w_4_19_1);
	full_adder (w_3_18_4, w_3_18_5, w_3_18_6, w_4_18_4, w_4_19_2);
	full_adder (w_3_19_1, w_3_19_2, w_3_19_3, w_4_19_3, w_4_20_1);
	full_adder (w_3_19_4, w_3_19_5, w_3_19_6, w_4_19_4, w_4_20_2);
	full_adder (w_3_20_1, w_3_20_2, w_3_20_3, w_4_20_3, w_4_21_1);
	full_adder (w_3_20_4, w_3_20_5, w_3_20_6, w_4_20_4, w_4_21_2);
	full_adder (w_3_21_1, w_3_21_2, w_3_21_3, w_4_21_3, w_4_22_1);
	full_adder (w_3_21_4, w_3_21_5, w_3_21_6, w_4_21_4, w_4_22_2);
	full_adder (w_3_22_1, w_3_22_2, w_3_22_3, w_4_22_3, w_4_23_1);
	full_adder (w_3_22_4, w_3_22_5, w_3_22_6, w_4_22_4, w_4_23_2);
	full_adder (w_3_23_1, w_3_23_2, w_3_23_3, w_4_23_3, w_4_24_1);
	full_adder (w_3_23_4, w_3_23_5, w_3_23_6, w_4_23_4, w_4_24_2);
	full_adder (w_3_24_1, w_3_24_2, w_3_24_3, w_4_24_3, w_4_25_1);
	full_adder (w_3_24_4, w_3_24_5, w_3_24_6, w_4_24_4, w_4_25_2);
	half_adder (w_3_24_7, w_3_24_8, w_4_24_5, w_4_25_3);
	full_adder (w_3_25_1, w_3_25_2, w_3_25_3, w_4_25_4, w_4_26_1);
	full_adder (w_3_25_4, w_3_25_5, w_3_25_6, w_4_25_5, w_4_26_2);
	half_adder (w_3_25_7, w_3_25_8, w_4_25_6, w_4_26_3);
	full_adder (w_3_26_1, w_3_26_2, w_3_26_3, w_4_26_4, w_4_27_1);
	full_adder (w_3_26_4, w_3_26_5, w_3_26_6, w_4_26_5, w_4_27_2);
	half_adder (w_3_26_7, w_3_26_8, w_4_26_6, w_4_27_3);
	full_adder (w_3_27_1, w_3_27_2, w_3_27_3, w_4_27_4, w_4_28_1);
	full_adder (w_3_27_4, w_3_27_5, w_3_27_6, w_4_27_5, w_4_28_2);
	full_adder (w_3_27_7, w_3_27_8, a27b0, w_4_27_6, w_4_28_3);
	full_adder (w_3_28_1, w_3_28_2, w_3_28_3, w_4_28_4, w_4_29_1);
	full_adder (w_3_28_4, w_3_28_5, w_3_28_6, w_4_28_5, w_4_29_2);
	full_adder (w_3_28_7, w_3_28_8, w_1_28_19, w_4_28_6, w_4_29_3);
	full_adder (w_3_29_1, w_3_29_2, w_3_29_3, w_4_29_4, w_4_30_1);
	full_adder (w_3_29_4, w_3_29_5, w_3_29_6, w_4_29_5, w_4_30_2);
	full_adder (w_3_29_7, w_3_29_8, w_2_29_13, w_4_29_6, w_4_30_3);
	full_adder (w_3_30_1, w_3_30_2, w_3_30_3, w_4_30_4, w_4_31_1);
	full_adder (w_3_30_4, w_3_30_5, w_3_30_6, w_4_30_5, w_4_31_2);
	full_adder (w_3_30_7, w_3_30_8, w_3_30_9, w_4_30_6, w_4_31_3);
	full_adder (w_3_31_1, w_3_31_2, w_3_31_3, w_4_31_4, w_4_32_1);
	full_adder (w_3_31_4, w_3_31_5, w_3_31_6, w_4_31_5, w_4_32_2);
	full_adder (w_3_31_7, w_3_31_8, w_3_31_9, w_4_31_6, w_4_32_3);
	full_adder (w_3_32_1, w_3_32_2, w_3_32_3, w_4_32_4, w_4_33_1);
	full_adder (w_3_32_4, w_3_32_5, w_3_32_6, w_4_32_5, w_4_33_2);
	full_adder (w_3_32_7, w_3_32_8, w_3_32_9, w_4_32_6, w_4_33_3);
	full_adder (w_3_33_1, w_3_33_2, w_3_33_3, w_4_33_4, w_4_34_1);
	full_adder (w_3_33_4, w_3_33_5, w_3_33_6, w_4_33_5, w_4_34_2);
	full_adder (w_3_33_7, w_3_33_8, w_3_33_9, w_4_33_6, w_4_34_3);
	full_adder (w_3_34_1, w_3_34_2, w_3_34_3, w_4_34_4, w_4_35_1);
	full_adder (w_3_34_4, w_3_34_5, w_3_34_6, w_4_34_5, w_4_35_2);
	full_adder (w_3_34_7, w_3_34_8, w_3_34_9, w_4_34_6, w_4_35_3);
	full_adder (w_3_35_1, w_3_35_2, w_3_35_3, w_4_35_4, w_4_36_1);
	full_adder (w_3_35_4, w_3_35_5, w_3_35_6, w_4_35_5, w_4_36_2);
	full_adder (w_3_35_7, w_3_35_8, w_3_35_9, w_4_35_6, w_4_36_3);
	full_adder (w_3_36_1, w_3_36_2, w_3_36_3, w_4_36_4, w_4_37_1);
	full_adder (w_3_36_4, w_3_36_5, w_3_36_6, w_4_36_5, w_4_37_2);
	full_adder (w_3_36_7, w_3_36_8, w_3_36_9, w_4_36_6, w_4_37_3);
	full_adder (w_3_37_1, w_3_37_2, w_3_37_3, w_4_37_4, w_4_38_1);
	full_adder (w_3_37_4, w_3_37_5, w_3_37_6, w_4_37_5, w_4_38_2);
	half_adder (w_3_37_7, w_3_37_8, w_4_37_6, w_4_38_3);
	full_adder (w_3_38_1, w_3_38_2, w_3_38_3, w_4_38_4, w_4_39_1);
	full_adder (w_3_38_4, w_3_38_5, w_3_38_6, w_4_38_5, w_4_39_2);
	half_adder (w_3_38_7, w_3_38_8, w_4_38_6, w_4_39_3);
	full_adder (w_3_39_1, w_3_39_2, w_3_39_3, w_4_39_4, w_4_40_1);
	full_adder (w_3_39_4, w_3_39_5, w_3_39_6, w_4_39_5, w_4_40_2);
	half_adder (w_3_39_7, w_3_39_8, w_4_39_6, w_4_40_3);
	full_adder (w_3_40_1, w_3_40_2, w_3_40_3, w_4_40_4, w_4_41_1);
	full_adder (w_3_40_4, w_3_40_5, w_3_40_6, w_4_40_5, w_4_41_2);
	half_adder (w_3_40_7, w_3_40_8, w_4_40_6, w_4_41_3);
	full_adder (w_3_41_1, w_3_41_2, w_3_41_3, w_4_41_4, w_4_42_1);
	full_adder (w_3_41_4, w_3_41_5, w_3_41_6, w_4_41_5, w_4_42_2);
	half_adder (w_3_41_7, w_3_41_8, w_4_41_6, w_4_42_3);
	full_adder (w_3_42_1, w_3_42_2, w_3_42_3, w_4_42_4, w_4_43_1);
	full_adder (w_3_42_4, w_3_42_5, w_3_42_6, w_4_42_5, w_4_43_2);
	half_adder (w_3_42_7, w_2_42_10, w_4_42_6, w_4_43_3);
	full_adder (w_3_43_1, w_3_43_2, w_3_43_3, w_4_43_4, w_4_44_1);
	full_adder (w_3_43_4, w_3_43_5, w_3_43_6, w_4_43_5, w_4_44_2);
	full_adder (w_3_44_1, w_3_44_2, w_3_44_3, w_4_44_3, w_4_45_1);
	full_adder (w_3_44_4, w_3_44_5, w_3_44_6, w_4_44_4, w_4_45_2);
	full_adder (w_3_45_1, w_3_45_2, w_3_45_3, w_4_45_3, w_4_46_1);
	full_adder (w_3_45_4, w_3_45_5, w_3_45_6, w_4_45_4, w_4_46_2);
	full_adder (w_3_46_1, w_3_46_2, w_3_46_3, w_4_46_3, w_4_47_1);
	full_adder (w_3_46_4, w_3_46_5, w_3_46_6, w_4_46_4, w_4_47_2);
	full_adder (w_3_47_1, w_3_47_2, w_3_47_3, w_4_47_3, w_4_48_1);
	full_adder (w_3_47_4, w_3_47_5, w_3_47_6, w_4_47_4, w_4_48_2);
	full_adder (w_3_48_1, w_3_48_2, w_3_48_3, w_4_48_3, w_4_49_1);
	full_adder (w_3_48_4, w_3_48_5, w_3_48_6, w_4_48_4, w_4_49_2);
	full_adder (w_3_49_1, w_3_49_2, w_3_49_3, w_4_49_3, w_4_50_1);
	full_adder (w_3_49_4, w_3_49_5, w_1_49_10, w_4_49_4, w_4_50_2);
	full_adder (w_3_50_1, w_3_50_2, w_3_50_3, w_4_50_3, w_4_51_1);
	half_adder (w_3_50_4, not_a31b19, w_4_50_4, w_4_51_2);
	full_adder (w_3_51_1, w_3_51_2, w_3_51_3, w_4_51_3, w_4_52_1);
	full_adder (w_3_52_1, w_3_52_2, w_3_52_3, w_4_52_2, w_4_53_1);
	full_adder (w_3_53_1, w_3_53_2, w_3_53_3, w_4_53_2, w_4_54_1);
	full_adder (w_3_54_1, w_3_54_2, w_3_54_3, w_4_54_2, w_4_55_1);
	full_adder (w_3_55_1, w_3_55_2, w_3_55_3, w_4_55_2, w_4_56_1);
	full_adder (w_3_56_1, w_3_56_2, w_2_56_4, w_4_56_2, w_4_57_1);
	full_adder (w_3_57_1, w_3_57_2, w_1_57_4, w_4_57_2, w_4_58_1);
	half_adder (w_3_58_1, w_3_58_2, w_4_58_2, w_4_59_1);
	half_adder (w_3_59_1, w_3_59_2, w_4_59_2, w_4_60_1);
	half_adder (w_3_60_1, w_3_60_2, w_4_60_2, w_4_61_1);
	half_adder (w_3_61_1, w_3_61_2, w_4_61_2, w_4_62_1);
	half_adder (w_3_62_1, w_3_62_2, w_4_62_2, w_4_63_1);
	half_adder (w_3_63_1, w_3_63_2, w_4_63_2, w_4_64_1);
	half_adder (w_4_5_1, w_4_5_2, w_5_5_1, w_5_6_1);
	half_adder (w_4_6_1, w_4_6_2, w_5_6_2, w_5_7_1);
	half_adder (w_4_7_1, w_4_7_2, w_5_7_2, w_5_8_1);
	half_adder (w_4_8_1, w_4_8_2, w_5_8_2, w_5_9_1);
	half_adder (w_4_9_1, w_4_9_2, w_5_9_2, w_5_10_1);
	full_adder (w_4_10_1, w_4_10_2, w_3_10_4, w_5_10_2, w_5_11_1);
	full_adder (w_4_11_1, w_4_11_2, w_3_11_4, w_5_11_2, w_5_12_1);
	full_adder (w_4_12_1, w_4_12_2, w_3_12_4, w_5_12_2, w_5_13_1);
	full_adder (w_4_13_1, w_4_13_2, w_3_13_4, w_5_13_2, w_5_14_1);
	full_adder (w_4_14_1, w_4_14_2, w_4_14_3, w_5_14_2, w_5_15_1);
	full_adder (w_4_15_1, w_4_15_2, w_4_15_3, w_5_15_2, w_5_16_1);
	full_adder (w_4_16_1, w_4_16_2, w_4_16_3, w_5_16_2, w_5_17_1);
	full_adder (w_4_17_1, w_4_17_2, w_4_17_3, w_5_17_2, w_5_18_1);
	full_adder (w_4_18_1, w_4_18_2, w_4_18_3, w_5_18_2, w_5_19_1);
	full_adder (w_4_19_1, w_4_19_2, w_4_19_3, w_5_19_2, w_5_20_1);
	full_adder (w_4_20_1, w_4_20_2, w_4_20_3, w_5_20_2, w_5_21_1);
	full_adder (w_4_21_1, w_4_21_2, w_4_21_3, w_5_21_2, w_5_22_1);
	half_adder (w_4_21_4, w_2_21_10, w_5_21_3, w_5_22_2);
	full_adder (w_4_22_1, w_4_22_2, w_4_22_3, w_5_22_3, w_5_23_1);
	half_adder (w_4_22_4, w_2_22_10, w_5_22_4, w_5_23_2);
	full_adder (w_4_23_1, w_4_23_2, w_4_23_3, w_5_23_3, w_5_24_1);
	half_adder (w_4_23_4, w_3_23_7, w_5_23_4, w_5_24_2);
	full_adder (w_4_24_1, w_4_24_2, w_4_24_3, w_5_24_3, w_5_25_1);
	half_adder (w_4_24_4, w_4_24_5, w_5_24_4, w_5_25_2);
	full_adder (w_4_25_1, w_4_25_2, w_4_25_3, w_5_25_3, w_5_26_1);
	full_adder (w_4_25_4, w_4_25_5, w_4_25_6, w_5_25_4, w_5_26_2);
	full_adder (w_4_26_1, w_4_26_2, w_4_26_3, w_5_26_3, w_5_27_1);
	full_adder (w_4_26_4, w_4_26_5, w_4_26_6, w_5_26_4, w_5_27_2);
	full_adder (w_4_27_1, w_4_27_2, w_4_27_3, w_5_27_3, w_5_28_1);
	full_adder (w_4_27_4, w_4_27_5, w_4_27_6, w_5_27_4, w_5_28_2);
	full_adder (w_4_28_1, w_4_28_2, w_4_28_3, w_5_28_3, w_5_29_1);
	full_adder (w_4_28_4, w_4_28_5, w_4_28_6, w_5_28_4, w_5_29_2);
	full_adder (w_4_29_1, w_4_29_2, w_4_29_3, w_5_29_3, w_5_30_1);
	full_adder (w_4_29_4, w_4_29_5, w_4_29_6, w_5_29_4, w_5_30_2);
	full_adder (w_4_30_1, w_4_30_2, w_4_30_3, w_5_30_3, w_5_31_1);
	full_adder (w_4_30_4, w_4_30_5, w_4_30_6, w_5_30_4, w_5_31_2);
	full_adder (w_4_31_1, w_4_31_2, w_4_31_3, w_5_31_3, w_5_32_1);
	full_adder (w_4_31_4, w_4_31_5, w_4_31_6, w_5_31_4, w_5_32_2);
	full_adder (w_4_32_1, w_4_32_2, w_4_32_3, w_5_32_3, w_5_33_1);
	full_adder (w_4_32_4, w_4_32_5, w_4_32_6, w_5_32_4, w_5_33_2);
	full_adder (w_4_33_1, w_4_33_2, w_4_33_3, w_5_33_3, w_5_34_1);
	full_adder (w_4_33_4, w_4_33_5, w_4_33_6, w_5_33_4, w_5_34_2);
	full_adder (w_4_34_1, w_4_34_2, w_4_34_3, w_5_34_3, w_5_35_1);
	full_adder (w_4_34_4, w_4_34_5, w_4_34_6, w_5_34_4, w_5_35_2);
	full_adder (w_4_35_1, w_4_35_2, w_4_35_3, w_5_35_3, w_5_36_1);
	full_adder (w_4_35_4, w_4_35_5, w_4_35_6, w_5_35_4, w_5_36_2);
	full_adder (w_4_36_1, w_4_36_2, w_4_36_3, w_5_36_3, w_5_37_1);
	full_adder (w_4_36_4, w_4_36_5, w_4_36_6, w_5_36_4, w_5_37_2);
	full_adder (w_4_37_1, w_4_37_2, w_4_37_3, w_5_37_3, w_5_38_1);
	full_adder (w_4_37_4, w_4_37_5, w_4_37_6, w_5_37_4, w_5_38_2);
	full_adder (w_4_38_1, w_4_38_2, w_4_38_3, w_5_38_3, w_5_39_1);
	full_adder (w_4_38_4, w_4_38_5, w_4_38_6, w_5_38_4, w_5_39_2);
	full_adder (w_4_39_1, w_4_39_2, w_4_39_3, w_5_39_3, w_5_40_1);
	full_adder (w_4_39_4, w_4_39_5, w_4_39_6, w_5_39_4, w_5_40_2);
	full_adder (w_4_40_1, w_4_40_2, w_4_40_3, w_5_40_3, w_5_41_1);
	full_adder (w_4_40_4, w_4_40_5, w_4_40_6, w_5_40_4, w_5_41_2);
	full_adder (w_4_41_1, w_4_41_2, w_4_41_3, w_5_41_3, w_5_42_1);
	full_adder (w_4_41_4, w_4_41_5, w_4_41_6, w_5_41_4, w_5_42_2);
	full_adder (w_4_42_1, w_4_42_2, w_4_42_3, w_5_42_3, w_5_43_1);
	full_adder (w_4_42_4, w_4_42_5, w_4_42_6, w_5_42_4, w_5_43_2);
	full_adder (w_4_43_1, w_4_43_2, w_4_43_3, w_5_43_3, w_5_44_1);
	full_adder (w_4_43_4, w_4_43_5, w_2_43_10, w_5_43_4, w_5_44_2);
	full_adder (w_4_44_1, w_4_44_2, w_4_44_3, w_5_44_3, w_5_45_1);
	half_adder (w_4_44_4, w_2_44_10, w_5_44_4, w_5_45_2);
	full_adder (w_4_45_1, w_4_45_2, w_4_45_3, w_5_45_3, w_5_46_1);
	full_adder (w_4_46_1, w_4_46_2, w_4_46_3, w_5_46_2, w_5_47_1);
	full_adder (w_4_47_1, w_4_47_2, w_4_47_3, w_5_47_2, w_5_48_1);
	full_adder (w_4_48_1, w_4_48_2, w_4_48_3, w_5_48_2, w_5_49_1);
	full_adder (w_4_49_1, w_4_49_2, w_4_49_3, w_5_49_2, w_5_50_1);
	full_adder (w_4_50_1, w_4_50_2, w_4_50_3, w_5_50_2, w_5_51_1);
	full_adder (w_4_51_1, w_4_51_2, w_4_51_3, w_5_51_2, w_5_52_1);
	full_adder (w_4_52_1, w_4_52_2, w_3_52_4, w_5_52_2, w_5_53_1);
	full_adder (w_4_53_1, w_4_53_2, w_3_53_4, w_5_53_2, w_5_54_1);
	full_adder (w_4_54_1, w_4_54_2, w_3_54_4, w_5_54_2, w_5_55_1);
	full_adder (w_4_55_1, w_4_55_2, w_2_55_4, w_5_55_2, w_5_56_1);
	half_adder (w_4_56_1, w_4_56_2, w_5_56_2, w_5_57_1);
	half_adder (w_4_57_1, w_4_57_2, w_5_57_2, w_5_58_1);
	half_adder (w_4_58_1, w_4_58_2, w_5_58_2, w_5_59_1);
	half_adder (w_4_59_1, w_4_59_2, w_5_59_2, w_5_60_1);
	half_adder (w_4_60_1, w_4_60_2, w_5_60_2, w_5_61_1);
	half_adder (w_4_61_1, w_4_61_2, w_5_61_2, w_5_62_1);
	half_adder (w_4_62_1, w_4_62_2, w_5_62_2, w_5_63_1);
	half_adder (w_4_63_1, w_4_63_2, w_5_63_2, w_5_64_1);
	half_adder (w_4_64_1, w_3_64_1, w_5_64_2, w_5_65_1);
	half_adder (w_5_6_1, w_5_6_2, w_6_6_1, w_6_7_1);
	half_adder (w_5_7_1, w_5_7_2, w_6_7_2, w_6_8_1);
	half_adder (w_5_8_1, w_5_8_2, w_6_8_2, w_6_9_1);
	half_adder (w_5_9_1, w_5_9_2, w_6_9_2, w_6_10_1);
	half_adder (w_5_10_1, w_5_10_2, w_6_10_2, w_6_11_1);
	half_adder (w_5_11_1, w_5_11_2, w_6_11_2, w_6_12_1);
	half_adder (w_5_12_1, w_5_12_2, w_6_12_2, w_6_13_1);
	half_adder (w_5_13_1, w_5_13_2, w_6_13_2, w_6_14_1);
	half_adder (w_5_14_1, w_5_14_2, w_6_14_2, w_6_15_1);
	full_adder (w_5_15_1, w_5_15_2, w_4_15_4, w_6_15_2, w_6_16_1);
	full_adder (w_5_16_1, w_5_16_2, w_4_16_4, w_6_16_2, w_6_17_1);
	full_adder (w_5_17_1, w_5_17_2, w_4_17_4, w_6_17_2, w_6_18_1);
	full_adder (w_5_18_1, w_5_18_2, w_4_18_4, w_6_18_2, w_6_19_1);
	full_adder (w_5_19_1, w_5_19_2, w_4_19_4, w_6_19_2, w_6_20_1);
	full_adder (w_5_20_1, w_5_20_2, w_4_20_4, w_6_20_2, w_6_21_1);
	full_adder (w_5_21_1, w_5_21_2, w_5_21_3, w_6_21_2, w_6_22_1);
	full_adder (w_5_22_1, w_5_22_2, w_5_22_3, w_6_22_2, w_6_23_1);
	full_adder (w_5_23_1, w_5_23_2, w_5_23_3, w_6_23_2, w_6_24_1);
	full_adder (w_5_24_1, w_5_24_2, w_5_24_3, w_6_24_2, w_6_25_1);
	full_adder (w_5_25_1, w_5_25_2, w_5_25_3, w_6_25_2, w_6_26_1);
	full_adder (w_5_26_1, w_5_26_2, w_5_26_3, w_6_26_2, w_6_27_1);
	full_adder (w_5_27_1, w_5_27_2, w_5_27_3, w_6_27_2, w_6_28_1);
	full_adder (w_5_28_1, w_5_28_2, w_5_28_3, w_6_28_2, w_6_29_1);
	full_adder (w_5_29_1, w_5_29_2, w_5_29_3, w_6_29_2, w_6_30_1);
	full_adder (w_5_30_1, w_5_30_2, w_5_30_3, w_6_30_2, w_6_31_1);
	full_adder (w_5_31_1, w_5_31_2, w_5_31_3, w_6_31_2, w_6_32_1);
	half_adder (w_5_31_4, w_3_31_10, w_6_31_3, w_6_32_2);
	full_adder (w_5_32_1, w_5_32_2, w_5_32_3, w_6_32_3, w_6_33_1);
	half_adder (w_5_32_4, w_3_32_10, w_6_32_4, w_6_33_2);
	full_adder (w_5_33_1, w_5_33_2, w_5_33_3, w_6_33_3, w_6_34_1);
	half_adder (w_5_33_4, w_3_33_10, w_6_33_4, w_6_34_2);
	full_adder (w_5_34_1, w_5_34_2, w_5_34_3, w_6_34_3, w_6_35_1);
	half_adder (w_5_34_4, w_3_34_10, w_6_34_4, w_6_35_2);
	full_adder (w_5_35_1, w_5_35_2, w_5_35_3, w_6_35_3, w_6_36_1);
	half_adder (w_5_35_4, w_3_35_10, w_6_35_4, w_6_36_2);
	full_adder (w_5_36_1, w_5_36_2, w_5_36_3, w_6_36_3, w_6_37_1);
	half_adder (w_5_36_4, w_2_36_13, w_6_36_4, w_6_37_2);
	full_adder (w_5_37_1, w_5_37_2, w_5_37_3, w_6_37_3, w_6_38_1);
	full_adder (w_5_38_1, w_5_38_2, w_5_38_3, w_6_38_2, w_6_39_1);
	full_adder (w_5_39_1, w_5_39_2, w_5_39_3, w_6_39_2, w_6_40_1);
	full_adder (w_5_40_1, w_5_40_2, w_5_40_3, w_6_40_2, w_6_41_1);
	full_adder (w_5_41_1, w_5_41_2, w_5_41_3, w_6_41_2, w_6_42_1);
	full_adder (w_5_42_1, w_5_42_2, w_5_42_3, w_6_42_2, w_6_43_1);
	full_adder (w_5_43_1, w_5_43_2, w_5_43_3, w_6_43_2, w_6_44_1);
	full_adder (w_5_44_1, w_5_44_2, w_5_44_3, w_6_44_2, w_6_45_1);
	full_adder (w_5_45_1, w_5_45_2, w_5_45_3, w_6_45_2, w_6_46_1);
	full_adder (w_5_46_1, w_5_46_2, w_4_46_4, w_6_46_2, w_6_47_1);
	full_adder (w_5_47_1, w_5_47_2, w_4_47_4, w_6_47_2, w_6_48_1);
	full_adder (w_5_48_1, w_5_48_2, w_4_48_4, w_6_48_2, w_6_49_1);
	full_adder (w_5_49_1, w_5_49_2, w_4_49_4, w_6_49_2, w_6_50_1);
	full_adder (w_5_50_1, w_5_50_2, w_4_50_4, w_6_50_2, w_6_51_1);
	full_adder (w_5_51_1, w_5_51_2, w_3_51_4, w_6_51_2, w_6_52_1);
	half_adder (w_5_52_1, w_5_52_2, w_6_52_2, w_6_53_1);
	half_adder (w_5_53_1, w_5_53_2, w_6_53_2, w_6_54_1);
	half_adder (w_5_54_1, w_5_54_2, w_6_54_2, w_6_55_1);
	half_adder (w_5_55_1, w_5_55_2, w_6_55_2, w_6_56_1);
	half_adder (w_5_56_1, w_5_56_2, w_6_56_2, w_6_57_1);
	half_adder (w_5_57_1, w_5_57_2, w_6_57_2, w_6_58_1);
	half_adder (w_5_58_1, w_5_58_2, w_6_58_2, w_6_59_1);
	half_adder (w_5_59_1, w_5_59_2, w_6_59_2, w_6_60_1);
	half_adder (w_5_60_1, w_5_60_2, w_6_60_2, w_6_61_1);
	half_adder (w_5_61_1, w_5_61_2, w_6_61_2, w_6_62_1);
	half_adder (w_5_62_1, w_5_62_2, w_6_62_2, w_6_63_1);
	half_adder (w_5_63_1, w_5_63_2, w_6_63_2, w_6_64_1);
	half_adder (w_5_64_1, w_5_64_2, w_6_64_2, w_6_65_1);
	half_adder (w_6_7_1, w_6_7_2, w_7_7_1, w_7_8_1);
	half_adder (w_6_8_1, w_6_8_2, w_7_8_2, w_7_9_1);
	half_adder (w_6_9_1, w_6_9_2, w_7_9_2, w_7_10_1);
	half_adder (w_6_10_1, w_6_10_2, w_7_10_2, w_7_11_1);
	half_adder (w_6_11_1, w_6_11_2, w_7_11_2, w_7_12_1);
	half_adder (w_6_12_1, w_6_12_2, w_7_12_2, w_7_13_1);
	half_adder (w_6_13_1, w_6_13_2, w_7_13_2, w_7_14_1);
	half_adder (w_6_14_1, w_6_14_2, w_7_14_2, w_7_15_1);
	half_adder (w_6_15_1, w_6_15_2, w_7_15_2, w_7_16_1);
	half_adder (w_6_16_1, w_6_16_2, w_7_16_2, w_7_17_1);
	half_adder (w_6_17_1, w_6_17_2, w_7_17_2, w_7_18_1);
	half_adder (w_6_18_1, w_6_18_2, w_7_18_2, w_7_19_1);
	half_adder (w_6_19_1, w_6_19_2, w_7_19_2, w_7_20_1);
	half_adder (w_6_20_1, w_6_20_2, w_7_20_2, w_7_21_1);
	half_adder (w_6_21_1, w_6_21_2, w_7_21_2, w_7_22_1);
	full_adder (w_6_22_1, w_6_22_2, w_5_22_4, w_7_22_2, w_7_23_1);
	full_adder (w_6_23_1, w_6_23_2, w_5_23_4, w_7_23_2, w_7_24_1);
	full_adder (w_6_24_1, w_6_24_2, w_5_24_4, w_7_24_2, w_7_25_1);
	full_adder (w_6_25_1, w_6_25_2, w_5_25_4, w_7_25_2, w_7_26_1);
	full_adder (w_6_26_1, w_6_26_2, w_5_26_4, w_7_26_2, w_7_27_1);
	full_adder (w_6_27_1, w_6_27_2, w_5_27_4, w_7_27_2, w_7_28_1);
	full_adder (w_6_28_1, w_6_28_2, w_5_28_4, w_7_28_2, w_7_29_1);
	full_adder (w_6_29_1, w_6_29_2, w_5_29_4, w_7_29_2, w_7_30_1);
	full_adder (w_6_30_1, w_6_30_2, w_5_30_4, w_7_30_2, w_7_31_1);
	full_adder (w_6_31_1, w_6_31_2, w_6_31_3, w_7_31_2, w_7_32_1);
	full_adder (w_6_32_1, w_6_32_2, w_6_32_3, w_7_32_2, w_7_33_1);
	full_adder (w_6_33_1, w_6_33_2, w_6_33_3, w_7_33_2, w_7_34_1);
	full_adder (w_6_34_1, w_6_34_2, w_6_34_3, w_7_34_2, w_7_35_1);
	full_adder (w_6_35_1, w_6_35_2, w_6_35_3, w_7_35_2, w_7_36_1);
	full_adder (w_6_36_1, w_6_36_2, w_6_36_3, w_7_36_2, w_7_37_1);
	full_adder (w_6_37_1, w_6_37_2, w_6_37_3, w_7_37_2, w_7_38_1);
	full_adder (w_6_38_1, w_6_38_2, w_5_38_4, w_7_38_2, w_7_39_1);
	full_adder (w_6_39_1, w_6_39_2, w_5_39_4, w_7_39_2, w_7_40_1);
	full_adder (w_6_40_1, w_6_40_2, w_5_40_4, w_7_40_2, w_7_41_1);
	full_adder (w_6_41_1, w_6_41_2, w_5_41_4, w_7_41_2, w_7_42_1);
	full_adder (w_6_42_1, w_6_42_2, w_5_42_4, w_7_42_2, w_7_43_1);
	full_adder (w_6_43_1, w_6_43_2, w_5_43_4, w_7_43_2, w_7_44_1);
	full_adder (w_6_44_1, w_6_44_2, w_5_44_4, w_7_44_2, w_7_45_1);
	full_adder (w_6_45_1, w_6_45_2, w_4_45_4, w_7_45_2, w_7_46_1);
	half_adder (w_6_46_1, w_6_46_2, w_7_46_2, w_7_47_1);
	half_adder (w_6_47_1, w_6_47_2, w_7_47_2, w_7_48_1);
	half_adder (w_6_48_1, w_6_48_2, w_7_48_2, w_7_49_1);
	half_adder (w_6_49_1, w_6_49_2, w_7_49_2, w_7_50_1);
	half_adder (w_6_50_1, w_6_50_2, w_7_50_2, w_7_51_1);
	half_adder (w_6_51_1, w_6_51_2, w_7_51_2, w_7_52_1);
	half_adder (w_6_52_1, w_6_52_2, w_7_52_2, w_7_53_1);
	half_adder (w_6_53_1, w_6_53_2, w_7_53_2, w_7_54_1);
	half_adder (w_6_54_1, w_6_54_2, w_7_54_2, w_7_55_1);
	half_adder (w_6_55_1, w_6_55_2, w_7_55_2, w_7_56_1);
	half_adder (w_6_56_1, w_6_56_2, w_7_56_2, w_7_57_1);
	half_adder (w_6_57_1, w_6_57_2, w_7_57_2, w_7_58_1);
	half_adder (w_6_58_1, w_6_58_2, w_7_58_2, w_7_59_1);
	half_adder (w_6_59_1, w_6_59_2, w_7_59_2, w_7_60_1);
	half_adder (w_6_60_1, w_6_60_2, w_7_60_2, w_7_61_1);
	half_adder (w_6_61_1, w_6_61_2, w_7_61_2, w_7_62_1);
	half_adder (w_6_62_1, w_6_62_2, w_7_62_2, w_7_63_1);
	half_adder (w_6_63_1, w_6_63_2, w_7_63_2, w_7_64_1);
	half_adder (w_6_64_1, w_6_64_2, w_7_64_2, w_7_65_1);
	half_adder (w_6_65_1, w_5_65_1, w_7_65_2, w_7_66_1);
	half_adder (w_7_8_1, w_7_8_2, w_8_8_1, w_8_9_1);
	half_adder (w_7_9_1, w_7_9_2, w_8_9_2, w_8_10_1);
	half_adder (w_7_10_1, w_7_10_2, w_8_10_2, w_8_11_1);
	half_adder (w_7_11_1, w_7_11_2, w_8_11_2, w_8_12_1);
	half_adder (w_7_12_1, w_7_12_2, w_8_12_2, w_8_13_1);
	half_adder (w_7_13_1, w_7_13_2, w_8_13_2, w_8_14_1);
	half_adder (w_7_14_1, w_7_14_2, w_8_14_2, w_8_15_1);
	half_adder (w_7_15_1, w_7_15_2, w_8_15_2, w_8_16_1);
	half_adder (w_7_16_1, w_7_16_2, w_8_16_2, w_8_17_1);
	half_adder (w_7_17_1, w_7_17_2, w_8_17_2, w_8_18_1);
	half_adder (w_7_18_1, w_7_18_2, w_8_18_2, w_8_19_1);
	half_adder (w_7_19_1, w_7_19_2, w_8_19_2, w_8_20_1);
	half_adder (w_7_20_1, w_7_20_2, w_8_20_2, w_8_21_1);
	half_adder (w_7_21_1, w_7_21_2, w_8_21_2, w_8_22_1);
	half_adder (w_7_22_1, w_7_22_2, w_8_22_2, w_8_23_1);
	half_adder (w_7_23_1, w_7_23_2, w_8_23_2, w_8_24_1);
	half_adder (w_7_24_1, w_7_24_2, w_8_24_2, w_8_25_1);
	half_adder (w_7_25_1, w_7_25_2, w_8_25_2, w_8_26_1);
	half_adder (w_7_26_1, w_7_26_2, w_8_26_2, w_8_27_1);
	half_adder (w_7_27_1, w_7_27_2, w_8_27_2, w_8_28_1);
	half_adder (w_7_28_1, w_7_28_2, w_8_28_2, w_8_29_1);
	half_adder (w_7_29_1, w_7_29_2, w_8_29_2, w_8_30_1);
	half_adder (w_7_30_1, w_7_30_2, w_8_30_2, w_8_31_1);
	half_adder (w_7_31_1, w_7_31_2, w_8_31_2, w_8_32_1);
	full_adder (w_7_32_1, w_7_32_2, w_6_32_4, w_8_32_2, w_8_33_1);
	full_adder (w_7_33_1, w_7_33_2, w_6_33_4, w_8_33_2, w_8_34_1);
	full_adder (w_7_34_1, w_7_34_2, w_6_34_4, w_8_34_2, w_8_35_1);
	full_adder (w_7_35_1, w_7_35_2, w_6_35_4, w_8_35_2, w_8_36_1);
	full_adder (w_7_36_1, w_7_36_2, w_6_36_4, w_8_36_2, w_8_37_1);
	full_adder (w_7_37_1, w_7_37_2, w_5_37_4, w_8_37_2, w_8_38_1);
	half_adder (w_7_38_1, w_7_38_2, w_8_38_2, w_8_39_1);
	half_adder (w_7_39_1, w_7_39_2, w_8_39_2, w_8_40_1);
	half_adder (w_7_40_1, w_7_40_2, w_8_40_2, w_8_41_1);
	half_adder (w_7_41_1, w_7_41_2, w_8_41_2, w_8_42_1);
	half_adder (w_7_42_1, w_7_42_2, w_8_42_2, w_8_43_1);
	half_adder (w_7_43_1, w_7_43_2, w_8_43_2, w_8_44_1);
	half_adder (w_7_44_1, w_7_44_2, w_8_44_2, w_8_45_1);
	half_adder (w_7_45_1, w_7_45_2, w_8_45_2, w_8_46_1);
	half_adder (w_7_46_1, w_7_46_2, w_8_46_2, w_8_47_1);
	half_adder (w_7_47_1, w_7_47_2, w_8_47_2, w_8_48_1);
	half_adder (w_7_48_1, w_7_48_2, w_8_48_2, w_8_49_1);
	half_adder (w_7_49_1, w_7_49_2, w_8_49_2, w_8_50_1);
	half_adder (w_7_50_1, w_7_50_2, w_8_50_2, w_8_51_1);
	half_adder (w_7_51_1, w_7_51_2, w_8_51_2, w_8_52_1);
	half_adder (w_7_52_1, w_7_52_2, w_8_52_2, w_8_53_1);
	half_adder (w_7_53_1, w_7_53_2, w_8_53_2, w_8_54_1);
	half_adder (w_7_54_1, w_7_54_2, w_8_54_2, w_8_55_1);
	half_adder (w_7_55_1, w_7_55_2, w_8_55_2, w_8_56_1);
	half_adder (w_7_56_1, w_7_56_2, w_8_56_2, w_8_57_1);
	half_adder (w_7_57_1, w_7_57_2, w_8_57_2, w_8_58_1);
	half_adder (w_7_58_1, w_7_58_2, w_8_58_2, w_8_59_1);
	half_adder (w_7_59_1, w_7_59_2, w_8_59_2, w_8_60_1);
	half_adder (w_7_60_1, w_7_60_2, w_8_60_2, w_8_61_1);
	half_adder (w_7_61_1, w_7_61_2, w_8_61_2, w_8_62_1);
	half_adder (w_7_62_1, w_7_62_2, w_8_62_2, w_8_63_1);
	half_adder (w_7_63_1, w_7_63_2, w_8_63_2, w_8_64_1);
	half_adder (w_7_64_1, w_7_64_2, w_8_64_2, w_8_65_1);
	half_adder (w_7_65_1, w_7_65_2, w_8_65_2, w_8_66_1);
	assign result1[0]=a0b0;
	assign result2[0]=0;
	assign result1[1]=w_1_1_1;
	assign result2[1]=0;
	assign result1[2]=w_2_2_1;
	assign result2[2]=0;
	assign result1[3]=w_3_3_1;
	assign result2[3]=0;
	assign result1[4]=w_4_4_1;
	assign result2[4]=0;
	assign result1[5]=w_5_5_1;
	assign result2[5]=0;
	assign result1[6]=w_6_6_1;
	assign result2[6]=0;
	assign result1[7]=w_7_7_1;
	assign result2[7]=0;
	assign result1[8]=w_8_8_1;
	assign result2[8]=0;
	assign result1[9]=w_8_9_1;
	assign result2[9]=w_8_9_2;
	assign result1[10]=w_8_10_1;
	assign result2[10]=w_8_10_2;
	assign result1[11]=w_8_11_1;
	assign result2[11]=w_8_11_2;
	assign result1[12]=w_8_12_1;
	assign result2[12]=w_8_12_2;
	assign result1[13]=w_8_13_1;
	assign result2[13]=w_8_13_2;
	assign result1[14]=w_8_14_1;
	assign result2[14]=w_8_14_2;
	assign result1[15]=w_8_15_1;
	assign result2[15]=w_8_15_2;
	assign result1[16]=w_8_16_1;
	assign result2[16]=w_8_16_2;
	assign result1[17]=w_8_17_1;
	assign result2[17]=w_8_17_2;
	assign result1[18]=w_8_18_1;
	assign result2[18]=w_8_18_2;
	assign result1[19]=w_8_19_1;
	assign result2[19]=w_8_19_2;
	assign result1[20]=w_8_20_1;
	assign result2[20]=w_8_20_2;
	assign result1[21]=w_8_21_1;
	assign result2[21]=w_8_21_2;
	assign result1[22]=w_8_22_1;
	assign result2[22]=w_8_22_2;
	assign result1[23]=w_8_23_1;
	assign result2[23]=w_8_23_2;
	assign result1[24]=w_8_24_1;
	assign result2[24]=w_8_24_2;
	assign result1[25]=w_8_25_1;
	assign result2[25]=w_8_25_2;
	assign result1[26]=w_8_26_1;
	assign result2[26]=w_8_26_2;
	assign result1[27]=w_8_27_1;
	assign result2[27]=w_8_27_2;
	assign result1[28]=w_8_28_1;
	assign result2[28]=w_8_28_2;
	assign result1[29]=w_8_29_1;
	assign result2[29]=w_8_29_2;
	assign result1[30]=w_8_30_1;
	assign result2[30]=w_8_30_2;
	assign result1[31]=w_8_31_1;
	assign result2[31]=w_8_31_2;
	assign result1[32]=w_8_32_1;
	assign result2[32]=w_8_32_2;
	assign result1[33]=w_8_33_1;
	assign result2[33]=w_8_33_2;
	assign result1[34]=w_8_34_1;
	assign result2[34]=w_8_34_2;
	assign result1[35]=w_8_35_1;
	assign result2[35]=w_8_35_2;
	assign result1[36]=w_8_36_1;
	assign result2[36]=w_8_36_2;
	assign result1[37]=w_8_37_1;
	assign result2[37]=w_8_37_2;
	assign result1[38]=w_8_38_1;
	assign result2[38]=w_8_38_2;
	assign result1[39]=w_8_39_1;
	assign result2[39]=w_8_39_2;
	assign result1[40]=w_8_40_1;
	assign result2[40]=w_8_40_2;
	assign result1[41]=w_8_41_1;
	assign result2[41]=w_8_41_2;
	assign result1[42]=w_8_42_1;
	assign result2[42]=w_8_42_2;
	assign result1[43]=w_8_43_1;
	assign result2[43]=w_8_43_2;
	assign result1[44]=w_8_44_1;
	assign result2[44]=w_8_44_2;
	assign result1[45]=w_8_45_1;
	assign result2[45]=w_8_45_2;
	assign result1[46]=w_8_46_1;
	assign result2[46]=w_8_46_2;
	assign result1[47]=w_8_47_1;
	assign result2[47]=w_8_47_2;
	assign result1[48]=w_8_48_1;
	assign result2[48]=w_8_48_2;
	assign result1[49]=w_8_49_1;
	assign result2[49]=w_8_49_2;
	assign result1[50]=w_8_50_1;
	assign result2[50]=w_8_50_2;
	assign result1[51]=w_8_51_1;
	assign result2[51]=w_8_51_2;
	assign result1[52]=w_8_52_1;
	assign result2[52]=w_8_52_2;
	assign result1[53]=w_8_53_1;
	assign result2[53]=w_8_53_2;
	assign result1[54]=w_8_54_1;
	assign result2[54]=w_8_54_2;
	assign result1[55]=w_8_55_1;
	assign result2[55]=w_8_55_2;
	assign result1[56]=w_8_56_1;
	assign result2[56]=w_8_56_2;
	assign result1[57]=w_8_57_1;
	assign result2[57]=w_8_57_2;
	assign result1[58]=w_8_58_1;
	assign result2[58]=w_8_58_2;
	assign result1[59]=w_8_59_1;
	assign result2[59]=w_8_59_2;
	assign result1[60]=w_8_60_1;
	assign result2[60]=w_8_60_2;
	assign result1[61]=w_8_61_1;
	assign result2[61]=w_8_61_2;
	assign result1[62]=w_8_62_1;
	assign result2[62]=w_8_62_2;
	assign result1[63]=w_8_63_1;
	assign result2[63]=w_8_63_2;
	
	wire cout;
	wire [63:0] out_untruncated;

	cla_adder final_add(result1, result2, 0, out_untruncated, cout);
	assign out = out_untruncated[31:0];
	
endmodule